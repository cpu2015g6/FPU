library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity fputop is
  port(MCLK1: in std_logic;
       RS_TX: out std_logic);
  end fputop;

architecture VHDL of fputop is

component fmul
  port(clk: in std_logic;
       op1, op2:  in std_logic_vector(31 downto 0);
       ans:       out std_logic_vector(31 downto 0) := x"00000000"
       );
end component;

component u232c
  generic (wtime: std_logic_vector(15 downto 0) := x"1ADB");
  Port ( clk  : in  STD_LOGIC;
         data : in  STD_LOGIC_VECTOR (7 downto 0);
         go   : in  STD_LOGIC;
         busy : out STD_LOGIC;
         tx   : out STD_LOGIC);
end component;

  signal clk,iclk: std_logic;
  type rom_t is array(0 to 2252) of std_logic_vector(31 downto 0);
  constant rom: rom_t := ("01011001011110100011000000100001",
"01000101101111001100000111000100",
"01011111101110000111100010110110",
"10111111111101111000000101011001",
"01101000100101010101000101111010",
"11101001000100000101110100001111",
"01001010110010110110101101101001",
"01001011100101111001010111101000",
"01010110111100001110011011110010",
"10011100100011101010001000001100",
"01001011001100111110111010101001",
"10101000010010001000000010001110",
"10111100001000000000101111010100",
"11010010011101001000101000000001",
"01001111000110001110000110001101",
"10011100110100111110001000000000",
"10111100100001000111011000001011",
"00011001110110110100010001110111",
"11001001000101111110000100110100",
"11100101100010011011110000111101",
"01101111001000110110111001100101",
"10101011010001100111111000000001",
"11001000010010110011010110101010",
"00110100000111011000111110000111",
"10110000111000001000011100100100",
"10110011110001110000011101011110",
"00100101001011101000111110000011",
"00110001010110100000010101100000",
"11001000010100011000010010001101",
"10111010001100100110111101000110",
"01010000001010111000000000010001",
"00011101101100011011100000001011",
"00101110011011100001110110101110",
"10011111011110001010110010010001",
"00100010111000111001011000011100",
"10000010110111010001001011010101",
"11010110101010101001110101111011",
"11100001011001000001010100000100",
"01111000100110000000001001000011",
"01000111100010100010101110111011",
"00110111010010001110111010010101",
"00111111010110001110010111011110",
"10110111111011011101100110110100",
"11100011011000000010000111101111",
"01011011110100000011111000000101",
"10110101111010101010101010011010",
"11111000001001001100011111111010",
"01101110100101110000110010011010",
"10011100001111100010100001011111",
"01101100001000110000101001000111",
"11001000111100100011011010101110",
"11001101100001110001111101001011",
"10001011001010010100010101101100",
"00011001001100101011000010011010",
"11000010011100100011010000000001",
"10111010111010000111101010101111",
"00111101110110111111001100110011",
"01010111101100111110000001100011",
"10101110011001111001101100010011",
"11000110101000101011110001110000",
"01100000111000101100011001010011",
"00001111001010110110110101000100",
"00110000100101111101101101000100",
"11110110100011001101100101111100",
"10111000111110111011010100100111",
"01110000000010100111110011101000",
"11100000001100000001110001110100",
"11010111011110001101110101110101",
"01111000001010110011001111101001",
"11111111011001001001111010110111",
"10000001000000111001011110111010",
"01000000111010110000100101101111",
"11101000100010111100101111001010",
"10001100111010111001000010001100",
"00110110000000001010001100000010",
"10011100000101101111110111010000",
"11010111001110101110011110100011",
"00110011110111000111101000010001",
"11000010100111100111101110110011",
"10110110100110010011010101011011",
"00111001101111011011000111101100",
"01101111100101001110101010000011",
"00111110001000011110111000001111",
"01101110001111000110001111101110",
"10101001111111100100110000001111",
"01101101001101100001011101001101",
"11010111101101001110000100111000",
"11000100101011101111010011000010",
"10100000101111010011001011010110",
"00100110000000010100110101110001",
"10101010001001000100111011110110",
"11010010101111000001110010010000",
"00111101011100010111100010100011",
"00000010010011010011101011110010",
"01000010000010110100100110110100",
"00000100110111110101010000101111",
"10011001010001100011000101010111",
"01001100010010011001001100000001",
"10100110000111000000111010001100",
"01010100001001101010100001011110",
"10000111001110100110010011100110",
"10011011111100101011000000001000",
"11110100011100000111110000110011",
"00001100011111010110000111001001",
"11000001011011100000011010011010",
"10101101001110101001010010011111",
"11001010011001011100001001001101",
"00111000001001110111010010001111",
"11011010000000101111000111101110",
"10110010111001110010010101101101",
"01001101011011000111011011100101",
"00000011101101111101010111000010",
"01100100001111011101001010001001",
"00101000100010000101000000000000",
"11101011011110000011011101101111",
"11001010011111000000000011100110",
"01110110011101000101011101110000",
"11010110111110010110001010101111",
"01011110010101101100111101111111",
"11110101110100010100001010100001",
"00101000101111001001000111001100",
"10011100101101110000001011011010",
"10000110000001101100111001010011",
"00111110100011010101001000010100",
"01011100011110101010110000100111",
"01011011100010100110000100110000",
"01110101001010100000110001101110",
"10001100101000111010100101100000",
"11000010010110010110110011011000",
"01010111000111111010101001000110",
"11000110100000001100111101111111",
"11011110001000001010110100011010",
"10100100110101111001111011111110",
"01011001100100110001110000011001",
"10111110111101111100111111101101",
"11110110010010100001111011110011",
"10001101110111111101111100100111",
"01000100101100001100000100100101",
"01101010010110101000101101001110",
"11001010001100101010010101000011",
"11110101000110001000000111110001",
"00101110000111111011110001001111",
"01111001111001110011110100000011",
"01101000100100000100100011111101",
"00100001000110110010101010100000",
"01101111000000001000111110010011",
"01010000100110111101100010101100",
"11101111110101110010110101011101",
"00110111001110101100100001000010",
"11100111100111001111111101001000",
"01000101000110101010011101101010",
"00001011011111011011000000110000",
"00010001000110010100000111100100",
"01010101101100000101010101110100",
"10100101100101010111101000010100",
"10111011110011011110101110100110",
"10011111011111001011011100010111",
"00111011100001000011100001100110",
"10011011100000101000011000010101",
"00101010100001001100011111111001",
"10100011101111001111100000111011",
"10001110110001000000011100110110",
"00010110110011100101101110011111",
"11000101001110110010011111101011",
"10011100100101101101110100011011",
"10000100010110011001011101011111",
"11110101010000011000000100011001",
"00111010001001000111100011011001",
"00001011100001011001001001011101",
"01110010010001011110001101101100",
"00111110010011101000000010010101",
"00101001100000001010101110101110",
"00101100011110101100001100000011",
"00010110011111000001001101011000",
"10110111111110000111001100110011",
"11111100011101101100100101100010",
"01110100111011111000001000100101",
"00100010000011000100001101110110",
"00101100010100101001100000111001",
"00001110111001101100010101111100",
"00111101111101100001100110011001",
"11011100010101011001000101100000",
"11011010110011010100111100001101",
"01010001100101110001001001111010",
"10011000101000111100000010011111",
"10101010110000010100010011011111",
"00101101001100101111111010010101",
"10111001111101110111000010011011",
"10100111101011010000001001011110",
"00110110011011100011100111111110",
"01000001000101100010100010100011",
"00111000000010111011101111001100",
"01101101011010001100000011011100",
"00000100010011010001010011011011",
"00110010001110100111010101100110",
"11011110100010011111100111010000",
"10011100001001000101010001001000",
"00111011001100010010001011101100",
"00110101001110110111000110100010",
"01100001011011011001011111010110",
"01010111001011011111011101100000",
"01100010001001011101001101101000",
"00000111111010110000000101100001",
"00101010100110000011100111110101",
"11000001111000100111000111111101",
"10010111100101010000100000111010",
"00011010000000111101001110011111",
"01100101001110100100001110100001",
"00101001110110110111101110110100",
"01001111100111111011000111011100",
"00110001110001100111110100010101",
"00011110100001110001000101110000",
"00010000110100010111001011110110",
"10110110000111000001100110101010",
"01001011001111010010110011001111",
"11000001111001101011010010001010",
"10110010100101011010101100000110",
"10111100110001001100010001111101",
"00101111111001100001001110100001",
"00100111100100110110010111101111",
"11110000001011101011111101111001",
"11011000010010010011101100001110",
"11110011000111010110110011000101",
"10001111000111100010111011100000",
"01000010110000101000101111101010",
"10100111000111011010001010010100",
"00111001000000000011001010011101",
"10100000100111011110000011101001",
"00111100110011001101111001101000",
"00111100111100110011001111111101",
"00111010010000101010000010110111",
"10001110000001100001101100011110",
"01000000001000000010001000011100",
"10001110101001111100010110100010",
"10001011010111010100111011101011",
"11111000001101111011011011100110",
"01000100000111101101000110000111",
"00110100111111000111101101100011",
"00100111110001001011101110010100",
"00011101010000100000011101111000",
"00010111111100110111101100001101",
"01000100100110010000001100000110",
"00011101000100011000011101101011",
"01010011101101110011000111100110",
"11010101011011101101010001010111",
"11101001101010101110100001010111",
"10001110011011110000011011110100",
"01101000000011101010101100011011",
"10110111000001010011010110011110",
"00100101000000011101111100011000",
"10011100000100001111100101101101",
"10000001100100110001100000001110",
"00001011100100000000001100011011",
"11010110101010100100000001111010",
"10100010101111111000110010101011",
"10010110110010100110001010010110",
"10110000101000111101011101101001",
"00001000000000011000011100010001",
"10101000110110111000111001001111",
"10110000101000011101001001010010",
"00011010000010101100100011100001",
"11011000011001101000110111100110",
"00111100010010001110001101111101",
"11010101001101001110101110111100",
"00000000111000011110011010000100",
"01000101011111100010100000000001",
"00000110111000000100011000000100",
"01000010000010001000001000011001",
"01100001110110101111000000001111",
"01100100011010010111110110010111",
"10111000100001010011000010001010",
"01011110001101110001101101010110",
"11010111001111101000011111010111",
"00001110110110101111001010111111",
"01000100111001101111011001101111",
"00010100010001011000100011011100",
"00001101110110101101001110010010",
"01001111111101100111010111000111",
"00011110010100101010101111111011",
"10010101011101001001110111001000",
"10111001101101000101000001100010",
"00001111101011000100101111000000",
"11011010101001001001011100101011",
"10110010110000111011111101100110",
"01001101111110111011010001101000",
"11011000101110110100100000010011",
"01001110010101011000011000010110",
"11100111100111000011010100010000",
"10110000001100000111011000100110",
"01001011011101011011100111010001",
"10111100001010010110000100101000",
"00101001101011001101010100100111",
"01001111100010101111001011001110",
"00111001101110111001110110100111",
"11111011000011100110111010000111",
"00000101110011001101001110110110",
"11000001011000111110101110111100",
"01010101110000110100100101111101",
"00010110001100110110100001000011",
"00101100100010001101101111101011",
"10101101101111111000111000011000",
"11110101010101110001111011010100",
"01100011101000001111011101100111",
"11000011101011001010010011101011",
"10011111110101000011001011101011",
"00100100000011110001101011101001",
"11101011010010011110110010111100",
"00001001100110101110111110111000",
"10110101011101000110101011111100",
"01011001001001011110001010000111",
"00010100100101111111101110010001",
"00101110010001001111011101000001",
"10111110000101000111101000000100",
"10111101101111001101001010111111",
"00111100010110110000011110101100",
"11000011100010011010011001110110",
"11001111011111001000011001101010",
"01010011100001111100100000100010",
"11010100101011011111010110000111",
"10100000000111100101100010100000",
"00110101010101110011001110000101",
"00010101011101010111011101110101",
"01101110010100111101000000000011",
"01000100010010110001100011101001",
"00110011110000011110100111011010",
"10101001100100011111100100110010",
"10011101110111010010010001101110",
"00111110001010011111010011000011",
"11011011111001110011101101011001",
"11011010100110011000001101000010",
"10011001101001000000111000011000",
"01110010000100100001010111101001",
"11001100001110110011110000101000",
"01000001100011101001110001010100",
"11110111011011011000000111111000",
"11111001100001000100111100100001",
"10011011000111011101010001011100",
"10111100111110100010100101111000",
"00011000100110100011101011110011",
"10101011010011011111100101111011",
"10110001001000110111101111000000",
"00011101000000111000100101101011",
"11011011010010100111010111100010",
"01010110101101001001111110100010",
"11110010100011101101100100100010",
"00000000010001101001100011010100",
"11000001010100001001110110100010",
"10000010001000011101011001110110",
"00001000100001011101101000101101",
"11110000000100000101001110110010",
"10111001000101101110110011111000",
"11100111011111011101010110101010",
"10001010100001000100000000100100",
"00110010100000110010000111000101",
"10000101100000111011101111011111",
"11001110001010010011001111010111",
"00010100001011100010001101100111",
"10110111110010011011101010000100",
"01011010111010100100010000111101",
"11010011001110001001101001000010",
"10110001100111101110001111011111",
"10100010110011110011111101000111",
"00010101000000001010000110000111",
"11100100000111111101110011101001",
"00111110000101001011110001000001",
"11100010101110011100001010001011",
"11010100100010001000000010000101",
"00101011000001010000011010101010",
"11000000000011011101110010100110",
"00011011000101010101101001011100",
"01001100001111010011100010011001",
"00100111110111001100100101110110",
"11010110110000010111100010111101",
"10011000011101011101001010110111",
"00101111101110011100011111001100",
"01100110100111110000011010001110",
"00011001100110111100101101001110",
"01000000110000011000111010000101",
"00100000010000100000101000010011",
"11001110000110111010000011100101",
"10101110111010111110110000011011",
"00101001000001011110010100100010",
"00011000000110110000110111011100",
"00000001101000100011000111110111",
"10111010111010100100110100100011",
"00001101010000001000010100100001",
"10001000101100000011001110110011",
"10100111111001010101011010101010",
"01011000100101010111110011100111",
"11000001000001011110101101010110",
"10100100110100101011010110000001",
"00100100000011101110110111001101",
"10001001011010110100100011010001",
"10011010010110100101101011011011",
"01010100110000000010011110110100",
"10101111101000111110011000000010",
"10100010110110111100100010011001",
"10111101000110011110010110011001",
"00100000100001000010000000000001",
"10101111111100010000110001110011",
"01001111100010110100101010010100",
"11000000000000110010011111111011",
"00101000001000001100011101111100",
"11110011001001111100001110000111",
"11011011110100101011100111011101",
"10010111001101101011000101010100",
"11100000010111101111010100110001",
"00111000000111110001110011000010",
"01100001000111011000010010111110",
"10100000011000010000111000010111",
"11000010000010100111101001010110",
"11110101001000010011010111001011",
"00001011110001010110001111011101",
"11000001011110001001101010010000",
"11001000110111110100100101110110",
"01001000101111000110111000001100",
"11010010001001000101100111101111",
"01000110100001001000110010010000",
"00001010011001010010001011011101",
"00010001011011010100011110010100",
"10111101011101011101111101010000",
"11011101010111001110100000101001",
"01011011010101000010101011100011",
"10101100111010000011001010111101",
"10011110001001101011110000101000",
"00001011100101110011101110010000",
"00010001010011100111111110101111",
"01100000000011100110001100000110",
"00110001111001011011010101100111",
"11000000011011010101100000110111",
"11101010100001000010001001110010",
"01101011011101010000001011011000",
"00001010111001010011000010001001",
"01110011000111111101101111001001",
"00111110100011110001110111101010",
"00011011110100110110111100100010",
"01111011111000100001000011010111",
"01011000001110101011011000000101",
"11010110011011111011000010101111",
"10010101010101101100111111100011",
"00101100010010010010000001010111",
"00100011001010110010110010100011",
"11010101011010101010001001101011",
"10111001000111001110001101100111",
"00101000100000011010001110000000",
"00100010110010011110110111101010",
"00001011110011001000001110110101",
"00011110101010111111111011000010",
"01001111101011011011101101101110",
"00101110111010010111001000101100",
"11100011101110011111111011111011",
"11011010100100100011101000111011",
"01111110110101000111101101110100",
"10110110011000100111101101011100",
"00011001110101000100010001000011",
"10010000101110111100101010001100",
"00010000001101011001000111101100",
"01100110110011101110000111010010",
"00110111100100101011101110010110",
"10011111011101001111010001111000",
"10110101111010100011000101011111",
"00010101111000000001011010110011",
"10110100010100010011111000000110",
"01001110100001011000001011001011",
"11000011010110100100000001000001",
"10110001010100111101001011011101",
"10011011110001011011110000100000",
"00001101101000111001110011101101",
"00001011001011110101111110111101",
"11101110110100100001100100001000",
"10111010100011111110110110101111",
"10100100101111000100101001101000",
"00110000001110101110111110000111",
"10010101100010010111111000111100",
"11000001110000100011111110100011",
"01010001111101010000001010110110",
"11010100001110011110100011110110",
"00100000011110101000010110000001",
"01011100000100110001111101101011",
"00111101000011111111100101101000",
"11111010111010111011011110101101",
"01000001000000010010100110110001",
"11111100011011011101101111100011",
"01100010001100000101100111100001",
"10000100010010101001111010000011",
"10100111000010111001010000011101",
"00000110111000110100100011100000",
"01101010011101111101100111110000",
"00110001110111000000110011001110",
"00011010101100101100100101110111",
"11000011001010001000001111100111",
"10011110011010110110000010101001",
"10010101000111011000011010011101",
"00111111100110000100011011111000",
"10010101001110110110011100110001",
"01011100100110100110101011101001",
"00110100111000001101000011001000",
"01010010000001111001101101111011",
"11001100100011000011100110011110",
"00101111000100011000000000111101",
"10111100000111110110010111000001",
"10110011010111000001111011000001",
"01000001000101001000001100001111",
"10110100111111110110010011110000",
"11011001001001011011001011100110",
"00000011001111100111000110010001",
"10011100111101101000100010010001",
"10010111101110001100011001000011",
"11100111010110010100000010001001",
"00111111100111001100111010100011",
"10100110111100011000011110000001",
"00110111011001101010010011011000",
"10011110110110011001101101000100",
"01010010111111111110011000010000",
"11010110101101000010100011011000",
"11101010001101000001011010010111",
"10001011100101001111100110100001",
"11100100001000011011010000101110",
"00110000001111000011001110110001",
"10010011001100110011010001101011",
"01001000001010011011101100001010",
"10011011111011011010000100010010",
"10001001001111100011111000011001",
"01001001000111101000011011111110",
"10010010111010111001110101001001",
"01001100010111001111100010001111",
"00011000101010000000000001010110",
"00100101100100010000001101101000",
"11101101001110000100001010110010",
"01001110000101010111101111010101",
"11111011110101110010111111100110",
"10110101011011101011110001011110",
"10100111010110100111011100011100",
"00011101010010111011101101111100",
"11011110110000010001101111110101",
"10010100001101011010111011010110",
"00110011100010010000110010100111",
"11011100010100101111000111100101",
"00001111001100011110110101001011",
"10101100000100101001110011000111",
"11010111010110111010100001010110",
"11010101011111011100101101001111",
"01101101010110011100001111001111",
"10011110100111000101001001001101",
"11010000000100010100011000001110",
"00101111001100010110101011001001",
"11101000101110010100011001100100",
"10000101011010101100010000110110",
"00101110101010011110100001011000",
"11010011100000000100000000001011",
"11100111100010001110011111110110",
"01111011100010010010110001110110",
"11111100011111011010111111000010",
"10000000110000001101000000001011",
"00111101101111110001000111111011",
"10001111111100101011110101010110",
"01010000111010000100010001001001",
"10100001010111000011110001010101",
"00100110011001100000111110011000",
"11111110011011000100000101110100",
"11100101010101000101000100110010",
"01001110011111011000011110000010",
"10001010111001100010001110001011",
"10011001111000111110101011110010",
"00010000010100001110011111000001",
"01010101000010000011101110110000",
"00100101110111100101011110100111",
"10111100100100010010001110100110",
"11101000000010101110100100001011",
"01100101000111011000001010101110",
"11010110010110111101011010001000",
"01011000011111100111101011001110",
"11101111010110101000100001010000",
"11011001001111110100101011011001",
"00100011101001100001010111001100",
"10111101011110000011010110100101",
"11110010011011010011000101011101",
"00011000011010001011100111111000",
"11001011010101111010000100001011",
"01100100111110101011010000000101",
"00000101010010011101110111000101",
"00101010110001011011000010000110",
"11101101010101001100011011010000",
"10000100001100010001000101000111",
"00110010000100110010101111010010",
"01010110010000000111010111000101",
"10100110000110010101100000100111",
"10111100111001101001000101010001",
"01111110100101111101001011110101",
"10011000111110111101010101111011",
"11011000000101010101101001110010",
"10111100101000011110101101001000",
"10101011000111111111101010001001",
"00101000010010100101111100110000",
"00101001111100100100110111010100",
"00101100000110110111101010011110",
"00010110100100110010100100101110",
"10111100000011011111001011110011",
"11001010100110100101101101110111",
"01000111001010110010110110111011",
"11001111111001000011100100111100",
"00011000010100011101110110101111",
"10101000101110110001100001011011",
"10011100100000101110111011110111",
"00101111100101001101100100001010",
"10001100100110000100001001010001",
"11010101101011100011000100110001",
"10010110111000001001011100110011",
"00101101000110001101000111101101",
"00101111110111000110110010101111",
"10011110110101011000001110100001",
"10001111001101111101011111000100",
"01001001111101010111111000101011",
"11101101001001100100011111110101",
"11110111100111110111010011010001",
"00010101111011101100011011111101",
"11001101000111010101100100011101",
"10100011100100101100001100100111",
"00010111101101111011010010010100",
"01110110110001000100010110011010",
"01001111000011001101100000110011",
"00001111000101100010001101001001",
"00110101100110011101111110001111",
"00000101001101000111110001100110",
"01100101001011101011100010011001",
"11000100000101111000010110100111",
"11101001110011101101010000110100",
"01011010111110000001110011011011",
"00111101101111000010100000000110",
"01011001001101100101101111111011",
"11011100100100011010101110100111",
"00111011010000000000111111101000",
"11011000010110101001001110010101",
"01111110110101001100101100110101",
"00001010010000100001011011011101",
"01001001101000010101010011111111",
"11010111010111110110111111111011",
"11000101100110111011001001001110",
"01011101100001111110010001101101",
"00111100010111111111011111101000",
"01011001110001011010110100001101",
"01010110101011001111000100101011",
"00001111010111111000110010011100",
"01111011100010000000000000111100",
"01001011011011011000010111001111",
"10111111100111111000010111100100",
"10010101011010111010010001101111",
"00010101100100101101011001011111",
"11010011001001111100110001110101",
"00111110100011100001110011110011",
"11010010001110100100110011000101",
"11111001110011100010110011011011",
"00011100101111110000110111001010",
"11010111000110011101111010010010",
"10110001110000001000110010011111",
"01100101110111100011010001011111",
"11011000001001110010000101010110",
"11110000001000000100101100111100",
"10011001000000110001010110110111",
"01001001101001000010100000110001",
"11011110100111101100100000000110",
"00101100000110010011011000101010",
"11001011001111100000111001001000",
"00001000110100011111001001100011",
"11011101100001000000100010010011",
"10100110110110001001000000000110",
"01110010111011111010110100000010",
"10111001001101111110010000001011",
"11101100101011000010101000101101",
"11110111110001100000000011111110",
"10001000011101010100011101001111",
"01000000101111011011011000011010",
"10100101001101000101010100011001",
"11001100000100011001001110000010",
"00110001110011010001100000110111",
"10110001111011111100011111100001",
"01011101000100110110101011110111",
"11001111100010100001001111110110",
"11111000111111000101100110111111",
"10100000001001101010111000011100",
"01011001101001000100110111010010",
"10101101011100001010000001000011",
"11010110001010001110001111000011",
"01000100000111101011111101000001",
"00110011101011001110110001010110",
"00011101111001100110000111010110",
"00010010000110111001111001101011",
"11010111000111100100010111100001",
"01100001101111010010010111110101",
"11111001011010011110001000011101",
"10101110100101101001011111100101",
"11010100010000010010011101001011",
"01000011011000110011111101000010",
"10110001010101001001001001000010",
"01101101111001011101110110100100",
"11011111101111101101111011011111",
"10111010110010010000000100111001",
"01101100001001100100000100111010",
"11100111100000101000101000000010",
"10001100010011001110111101010111",
"01101011110101000110010001001000",
"10111000101010100000011001111011",
"11000001111111010100100000001011",
"01000110101110100100010010111010",
"11001001001110000100101001010111",
"01010000011100010101001100100101",
"10001000111110101110000010001010",
"10011001111011000111111011011101",
"11101011011111111110010011101101",
"01001011000110111010100000001011",
"11110111000110111001011110010101",
"10011111010111001100111101010110",
"00110000011001100010011011011110",
"10010000010001101000001111001110",
"10011110010011000000010010000011",
"01111101001100110100111101111110",
"11011100000011101110011010000001",
"01100000000100010011010001110110",
"10111111011110101111100010100011",
"11100000000011100101101001000011",
"00001110000110000101111100011100",
"10110011111111110111111010011110",
"10000010100110000001001000011010",
"00111100111110100101111100101000",
"10110001001110000000001110110010",
"10101110101100111111100000000010",
"00010011100111100001110001010000",
"10111101001011011001110110000001",
"10010001010101100111010011010010",
"10111010011000001110110011111111",
"01100100011111100101000100110101",
"11011111010111110111001001111111",
"01011000101110110010000101100011",
"10010111110110011000011101000011",
"10110001000111110000001000101100",
"11010111010101000111111111100110",
"01001000110001010000110101110011",
"11100000101000111001000110010110",
"00100110100100110000000111011100",
"01101110111101000111000110010010",
"01010110000011000101111011111101",
"10100000001011000111010101000100",
"11101101111110001100001101100110",
"01001110101001111001010100111100",
"11010001001100001011100011011000",
"11001110100110000110011000000001",
"01100000010100100110100001010101",
"11101000000001101001011011001110",
"00110110110011111000001000101100",
"11011111010110100011000011000001",
"10100101110000111111001110111110",
"01111111001111011010100000001011",
"11100101100100010010101110010100",
"11001100110001110000010011001001",
"10011010101000010010011000011001",
"00100111111110101000111101000001",
"10111111001100111001111011011011",
"00111001111011101110111101110000",
"10111001101001111010010110101111",
"11011011101001110000101111111100",
"10001000100101010110011100000111",
"00100100110000101111101001101000",
"10001011110101111101001100001001",
"11000100101010001001010101100010",
"00010001000011100010000001101110",
"10111010000110111010100011110001",
"10010100100011101011010001111011",
"00001111001011011000101011100111",
"01001011010111100011011010100111",
"10110110100000100101110010100011",
"11000010011000100101000001010100",
"10110101110000000000010010101110",
"00100010111000101101001000011001",
"10011001001010100010000110111000",
"10111110100000100111110101001110",
"01100101000110010111011011000011",
"11100100000111000111001011011010",
"10101010010101010011010011000001",
"01010101100000010000110010010111",
"11000000010101101111010000100011",
"00010011111110000101111101001001",
"00110111010011101111010111011100",
"00001011110010001100101100110101",
"01011010001100011100011111110101",
"01011101101000101011010110000111",
"01111000011000011111110100110010",
"11010010100111111111011001100010",
"00101111100000010010110001111000",
"11000010101000010110110111100001",
"10010100100110101010001100111011",
"01011010001111100100010000000111",
"10101111011001011101110001111011",
"00111111111010101110001101100110",
"11011010101011100011011000010001",
"11011011000111111101100000101011",
"10110000001011110100001010101000",
"11001101001101100010111100101101",
"00111101111110010111001101011111",
"00101010101011000011000111010011",
"11010101010001000001001101001011",
"11000000100000111110001100100000",
"10001100100100110000100100100111",
"01110110001111010001110110010110",
"11000011010110010011110110000000",
"01000011000110000011000110110001",
"11001011001000111011100001110100",
"11001110110000101010101010011001",
"11111010101001001110010011101100",
"00010100111100011011010101011100",
"11010000000110111011000001010011",
"10111101010011111111111000010101",
"01000110111100000001000010101001",
"11000100110000110000101110111101",
"10111101001011010010111000111111",
"11001100001111010010001000111010",
"01001001111111111110010010011000",
"11000001010010001110101101101000",
"10010010101011111110001001001100",
"00010100100010100000101010001000",
"01011101110100111001101011000000",
"11010010011000100110001111110011",
"11110000101110110010000100111011",
"11100111010101000001100101001111",
"01000000111100111110000011101111",
"11101000110010100000111001100010",
"10010011000110100111100110101110",
"11111001010000010001000100000011",
"01001100111010010000000000000000",
"01011011001001100111111111010010",
"00101010010001010111111101101110",
"01000110000000000111001100111110",
"11110110100000101010000110101000",
"00111110111000001010110011011111",
"11110101111001010100101101010011",
"11010001100100001000111100101011",
"00000101011100110101011011011100",
"10010111100010010110100011110010",
"11010111110101011011101011001111",
"11010110010001011110111101010101",
"01101110101001010100000010010010",
"10010111001110011101000001000101",
"11101111100101001011000101101110",
"01000111010101111101101001100001",
"01101000110101011100001001110001",
"00011011010011001101011001001101",
"01000100101010110000100111100011",
"00111010010001101011101010111000",
"10000111001101101110110001100110",
"10000010000011100000000001000010",
"10011011011011010101101110001111",
"10110110111111110001011100000100",
"00010010111011001000001110001010",
"11100001010001001001011001110010",
"10010011110110110010101110111110",
"00110101101010000100111001001011",
"11010010101110111101100010011101",
"10111000010010000011100011100010",
"01001011100100101110101011111000",
"10111101101110111000111110111110",
"01001011101111110110111101010101",
"11001010000011000100000111010000",
"10100010000001010101111010101010",
"11011011100011010011101101001110",
"00111110000100110010100000010010",
"01001011001000011110110010111100",
"11101010011010010000010101111110",
"11110110000100110110001111110000",
"10000101101101011101101111001011",
"01001101110101110000101101010011",
"10010100000110001100001110100011",
"10011010110001101010001101100111",
"01110101111101101011100000011101",
"11010001001111110110111111100001",
"10101110001111101111000011111111",
"01110011100111110010110100100010",
"11100010011011010111001010110000",
"00111111010111101001110001110111",
"01100101011111110111010110000010",
"01100101010111100010010000001001",
"11000001000011001011000011010000",
"01010110010001101110100111111001",
"11010111110110101010001010101101",
"11000000101011111110111101110111",
"11111110001101101010001011110100",
"01111111011110110000100001111000",
"11001100000011011010111001000111",
"01100011100011100000101001100010",
"11110000000111010011100011010101",
"01010111100011111000110011000111",
"10000111101010111000001000111000",
"10011111110000000101100000011100",
"10001110100101101111100111100001",
"01111000101001100010011111110001",
"11000111110000111111101100101100",
"01100110100000001110101100100110",
"00101000101011101111110100011010",
"01001111101100000011111010010011",
"01100000101010010000011100010001",
"00100001111001101010110011010001",
"01000011000110000100111001110100",
"01110101110011001010010111001011",
"00011110110111011001110101010100",
"01010101001100010010100011100101",
"10010111100000111100010101000110",
"01101000000100110010000100011011",
"11000000000101110111011010100011",
"01011010111101001101111100011111",
"01000100101000010101011001000010",
"01100000000110100101001011010101",
"01101101010100000101001101011100",
"10101011110100101100100000101110",
"11011001101010111000011101001000",
"10110110001101001110010101000110",
"11101110100110001101010010100100",
"01100101010101111111110011000111",
"11000001101100111011100000010100",
"00011111111101011010010010101011",
"10100010001011000111001011000101",
"11001000111011000001000010101000",
"01110000101111010100000000010110",
"11111010001011101000001101100100",
"11011000110100000110000100110010",
"10110110000010000100101010101010",
"01001111010111011110000011010010",
"11111010101010011010000011101100",
"10001001100011001111000110100101",
"01000100101110101100100000111110",
"00110101010111111011100111010100",
"01011100100100000101110001111011",
"01010010011111000101001010110011",
"01001011001010010011000100011111",
"10101110001100101010001110101001",
"10111001111011000010000010100011",
"01010100010101100100111000001010",
"10111010101010010110111001010010",
"11001111100011011101010111011111",
"11011010100111110001001011111101",
"10101001000011010101001100010111",
"01000100001011111010001000101110",
"10101010111010001010000110100100",
"11100011000010000010100001000101",
"01001110011101110111010011101110",
"10111101011110011001001111111110",
"01110001000001001111000100011100",
"11101111000000011001101101011111",
"11001010101001010110110010011101",
"11110000100100001111101110000011",
"01111011101110110101111100111101",
"00011001100111100100111010011010",
"01100000011100111011111100111001",
"00111010100101101011101011011100",
"01101111011100111111101100010101",
"10000101001110011001100100011100",
"10110101001100001110001001011110",
"01101000010000011100000101100010",
"11010001011111101010111101111000",
"11111010010000001100001010101101",
"00110010011001111110011011111011",
"11001101011110110001011000100100",
"11000000011000110111001110000111",
"10111110100000000000011101000001",
"10000100010101010010000111100101",
"00000011010101010010110111111001",
"10010100010100010010000000110001",
"01011100110011111011011111001010",
"10110001101010011010111100101011",
"11001101011000001011001101001101",
"01011010110111010110011111000111",
"11101000110000100101010111100000",
"00111011010100010010011100000000",
"00010010001101010110011101000000",
"00001110000101000011010011101110",
"10001100110010010000101101011011",
"01011100011110110000001100001000",
"10101001110001010010000010000100",
"11100001101101001001110000100100",
"00011101110110000100101000001001",
"11000000000110001001011111111010",
"01100110111101000101001101011000",
"10010001100000001011101010111000",
"10111000111101011011011111000000",
"11101100010111100010001001111111",
"10010001011100001100001100101110",
"00111110010100001110100110110011",
"10100011101001100010101001101110",
"11101111000011010001111101111011",
"01010011001101110011001110011011",
"11001011100010000010001010000011",
"01101001110101110100001010000110",
"11110101111001001111000010111000",
"00000111101011111000110010010000",
"11000011010001011101111101100010",
"10001011100001111011000001011001",
"00101011100110010011110011100001",
"00101010011001011100001000000100",
"00010110100010011000011110011000",
"00110100100010100101110110010001",
"11100000100100001101011000101001",
"11010101100111001001000011000100",
"11110010000100011001000011100001",
"00000000111111000010011101100001",
"10110011100011110110000100000010",
"10010010011011001110101010001111",
"11101011001001111100000000011100",
"00111110000110110011111011001101",
"01011010001101001101111110011000",
"10110111111011100111011111101000",
"11010010101010000111110010010111",
"01010110011101000110011001100001",
"01001010001011001101110011110010",
"01100001001001010000011110111000",
"11100000001011010011000111110100",
"10111001010000010011001110011110",
"01011010000000101011010110010101",
"01100011101001101111010110100010",
"01001110011010100101110011101111",
"01110010100110001101100100100010",
"10101110111110110011001100011000",
"11000101000101000010011000011000",
"00110100100100010101111011101011",
"11000110000100000100110101111001",
"00000011100000111011101110101100",
"10001010000101001000001011011101",
"11101110101010110111101111001001",
"10000101100110110111010000111000",
"00110100110100000100001110011001",
"00111101100010011110110000100001",
"01110101000100101001011111001011",
"01110011000111011111010011100101",
"10001000010000010001111011001010",
"01000001100101110001111001000000",
"10001010011000111111111111110110",
"01001011011101110110110011111010",
"11001001000001010101000101110111",
"11010101000000001101101001011010",
"00100000100101110100111110011110",
"10111011001101110100101000010111",
"10011100010110001010101101101001",
"10110000010010011110000111100011",
"10111011101101110010101110000101",
"00101100100100000111001011001011",
"00110101110000000101111110010000",
"01110110011110111001001110110001",
"01101100101111010000110010101110",
"10001000100001011100111011100011",
"11000100101011110101010001100010",
"00001101101101110100100100010001",
"11011111101010110010111111001000",
"11000100101010101001100100111011",
"01100100111001000010100001100100",
"10101011000111100011000111110110",
"10011011110101001001110101110110",
"00000111100000110110001010101101",
"01100110001100000001111011111010",
"10100110100000100011001011001111",
"11001101001100110010010101011111",
"00010011001111010100000011101000",
"00111011100110101100110100101011",
"00001111011001001110000101110001",
"00110010000101100110000011011100",
"10100001011000110100001011011100",
"10010100000001010111111100101001",
"01100110000100101001011100111110",
"10100100110110110001001111000001",
"11001011011110101110010101100100",
"01101010011001000011010001011011",
"10100100011001000000000110010100",
"11001111010010110100000000001001",
"11000000001110001001111100001010",
"10000010010010100001101101101001",
"00000011000100011100000101000010",
"10000010010000010110011100100110",
"11101111011011011010001010111111",
"00110010001100111000011101110010",
"11010010110110000100000111101011",
"10101010000110101101101011101010",
"00111101100000101101000010010101",
"10010011001101111111010111110000",
"10111101010011101100001001111001",
"00010001000101001001001110100110",
"01100001101100101100010000001110",
"00010000010111011101010100011011",
"00110010100110101110100000010000",
"10010010101001111111000010000101",
"11010001000011010111001010101001",
"00100100001110011001010101100010",
"01000000011110110001010101101001",
"00110111111100100111001110101001",
"00111000111011011100101110101110",
"11001111001011111110100001101001",
"00101111010000100110011000110000",
"10111111000001011001010001010111",
"00101001001011010110110100100100",
"10100010101011110001100001111111",
"10001100011011010011110001101000",
"10001010110010000101110010110001",
"01001110000110011001001100100001",
"10011001011100000110010100011010",
"01111101010110111111100101010001",
"00001010001110101000110011111000",
"01001000001000000100110001000110",
"01111011111111010100010101010110",
"10100010111101110011110010001001",
"11011111011101001001100111001010",
"10001001011110001101110000101010",
"11010010000000001010110100110001",
"00011011111110100010110011100011",
"10011111101110110011110100100010",
"00100011011010010110110111011100",
"10000011101010101011101011111110",
"00111100001110010000010111100100",
"00101001101110100010100101001011",
"00100110100001101000110000100000",
"11001100011010010100000111001010",
"10100110001010000001111110010100",
"00110011000110010010111111110010",
"00001001001110101000011000000110",
"11011001101111110001100111010101",
"10100011100010110011110011010001",
"01111100101101100101011001011110",
"00001111101111011110011000110001",
"01001101000001110100000110111000",
"01010010010010000100000100001110",
"11000011101111110000011000010100",
"11010110100101010110110101001011",
"11001011100111011000101010000010",
"11010011001101001011110101010000",
"01011111010111100111001111001000",
"11010010001101001011011001011110",
"11000100011010100011110111111010",
"01010111001001010101101001110010",
"00011110001010010101011111010000",
"01011101010010110000001100000110",
"00111100000001100100101010100010",
"01000101111111110100110001011100",
"10101111011100110101011100010001",
"10110101111100101010110001001111",
"11000000001111101011001101000011",
"01101000001011101111101111000110",
"11101001000000100101100101100101",
"11000001110100100000000001000010",
"00100111110100101000001010000111",
"10101010001011001010111101001001",
"10111000001000001101100010111111",
"11100010010000101110010010001110",
"01011010111101001110011110110110",
"10111111100011011110011110010100",
"10001001010100100011101001011101",
"00001001011010010001000010100011",
"11011011111100110011100110111000",
"00010010001110001011111101110100",
"10101110101011111000011101100011",
"11000001101011000001011010000101",
"11001011100111111001101010000011",
"01001101110101101001001110110100",
"01001000000111110100011110110001",
"00101110100000010101010101001001",
"00110111001000001111000001100001",
"10110100110001001110101001111111",
"10111111100011101101101100010010",
"00110100110110111100010100101010",
"10110011010001010111010111010110",
"11111111000100110000101010000010",
"01110010111000101101010110001010",
"01100001010101011110111100010000",
"10100101101100110101001100101001",
"11000111100101011101101110100111",
"00101111000001011000110110000110",
"00110010110110100101110111100010",
"00100010011000111101011011111101",
"01000101000100110001110101010110",
"01001000110110001111010011010101",
"01001110011110010101101011100110",
"10010100011110001000111101011000",
"00101011101001001101101010100000",
"10000000101000000001000000011010",
"01011010001001100010111111101001",
"01100100011000111110111001110001",
"01111111000100111111011101000110",
"11110001010101100101011001101001",
"00010111011110011010010111011111",
"11001001010100010000010011101101",
"11010111000010001000000011110001",
"10101111010010101010111001011110",
"01000110110110000010010101110000",
"10101110010111011011100011100000",
"01010010111011111000101111001100",
"11000001110011110111100010101101",
"11111000101000101101111011110101",
"00110111011001001100010010000001",
"11110000100100011000101110010111",
"01000110111010110001101011011011",
"01011111100011001000000100001101",
"01100111000000010000100100110100",
"00001011001100010101101110101101",
"01010110011111100010110011001011",
"00100010001100000001011111111110",
"00111010111000100001101100111101",
"00011100111100010101001100111100",
"00011000010101010010010100101000",
"00110100011010101111100100011011",
"00011111100001101101111011010111",
"00010100011101111001010111011011",
"01001110110100011000110100110101",
"10101000001110110001110111001101",
"10110111100110010010101010001011",
"11111011001010101010100110011001",
"10001011011101011011011000110001",
"01000111001000111100110111000101",
"11000010110110100111101010110010",
"00111101011110100110110010011011",
"11000000110101011011100010000010",
"00111011100011001001001010100001",
"01001110000101110010100011000101",
"01001010001001100000000111000000",
"00101101101000111010100111010010",
"10010010011111010101000001100110",
"10000000101000011111001000111011",
"11101000111110110111110100110001",
"00010101110101101101100011101110",
"10111111010100110000111111000010",
"00110010110010000010110000101011",
"01110100010110101001110110100011",
"01100111101010101111000011011111",
"01001010101001001101101001101111",
"10001000011010000001000000100111",
"10010011100101010111000001011011",
"00010011110111011100011001011000",
"01101100110001010011110111001010",
"01000001001010101101111100101001",
"00101010001111111010101001100101",
"01010101000100110000000110100011",
"00111111110111000010000000100011",
"00100011001010100010101001101000",
"11100000001111011011101011110000",
"11000011111111000011101100100010",
"01110010101110110000101101010110",
"01000110000111110100001000110011",
"01111001011010001011100011010001",
"01011011111101100001101100100001",
"00100111110011110110101011010000",
"01000100010001110110011010011111",
"10011100001010100000100001110011",
"01001111101010100010101100001011",
"10101100011000100000110001100110",
"11011111011001100001110000101100",
"10111100001001010101001010111110",
"01011100000101001001101010001000",
"10010001001110000101010001100001",
"11011111011010000000000110010000",
"00110001001001110000110110011000",
"00111111101001011011110010000000",
"11010111101101011110111000011001",
"11010111111010111001000011011000",
"00110110101000101001011110001111",
"00001101101010110111000101010101",
"00000100110110011100011001101111",
"11100111000100110000101100110011",
"00010101100101101011001110001110",
"10111101001011010001111101100101",
"11001010110011111101111100001111",
"00111000100001110010110100010101",
"11000011110110111000011001111000",
"10010111111011110010111010100101",
"11100000101101010111100001000100",
"00111001001010011000110001011000",
"00111000011010110110011001011101",
"00010101100110110000010100111110",
"00001110100011101000101111001100",
"00100101101110000111010010110001",
"11011000100101010111010011010010",
"10111110110101110110000000101110",
"11010111000100000111010000100000",
"10110000101101011000111001111111",
"01001000010011001110010100000101",
"01000110010011000100001000001101",
"11011110100110011101101101001010",
"11100101011101011000010011100011",
"00101011101011101101110101001110",
"10100111011001001111011011000110",
"10010011100111000110010110101001",
"10111010001000100011000110010010",
"10100101001010001010101000010101",
"00011111110101011011100010010100",
"10111101001101011010110101110001",
"01100110110100100100111000101001",
"11100100100101010011111110111111",
"10111111011001111100001011111100",
"01100111011111101001011010101001",
"11100111011001100111101111011011",
"10011000001101000010010100101000",
"10111000011100111100100001010011",
"00010001001010111000110000111100",
"00010111000011011010001110011101",
"11101010110100100101110100000011",
"11000010011010001100011101011010",
"10001010100010101011010000010001",
"11010000100000101100101111111110",
"00011011100011011011101111101110",
"10001101101000101001011110101101",
"01101001111100010110010010010100",
"10111000000110010101000010101011",
"01010000110000111011001010111110",
"01000111010111011011101010001110",
"01011000101010010111111111101010",
"00101110110111000101000100110111",
"00010011110000101001101001110100",
"00000011001001110111101001111000",
"11100110000100011100000001001001",
"01010010100101010001100011001000",
"11111001001010011100011000001101",
"10110101101110101101011000010011",
"10100011111111000110001110000001",
"00011010001110000011001101011010",
"01110100011111110010111101111111",
"10011010111110111010111010010000",
"11001111111110101110000110010011",
"01101101110011111001100110110110",
"10001001101101101110000000110101",
"10111000000101000100110100011001",
"01011011111000100101011110101011",
"00110100100010011111010101110010",
"01010000111100111111001111011010",
"11011000100001100101100011110011",
"00001010101010111000100011001100",
"10100011101101000000101001101001",
"10100101101001110011011101011100",
"10100100110011010110010100100100",
"00001011000001100010100101100101",
"11001010111000110000101011100111",
"11001111010001000000000111111000",
"01011010101011011101011000011000",
"11110101101101011110000100100000",
"00010110001001011000000001001111",
"11001100011010110010101010000101",
"10011111110111000110000010000100",
"10101100101010110000010100100101",
"00001101000100110011100011100110",
"11000100010001001110010011001011",
"11100011111011011100011100010001",
"01101000101101101110000011101011",
"10010111101010111000010001110010",
"00101100100111010100001101000001",
"10000100110100101011101010010010",
"11010001011010101010100001100101",
"00000100100111100010001110001100",
"10010110100100001111010010000100",
"01010011111000100010010110000100",
"00100000101001001001011010101110",
"00110101000100010110010100100100",
"00110110110010100001011011111110",
"00110010111011001001101011100001",
"00101010001110101100011101110110",
"01011111100101111010000000000111",
"00101101010011101110011100111101",
"01001101011101010001011101110110",
"10010001001111001010111001001110",
"00111011000000100000101101001101",
"10001100101111111011000110110000",
"10101110111110111010011110111111",
"11001011000000111101011101110101",
"00111010100000011001101010100100",
"01011000000000111101001100011011",
"10100010010011111001110100111111",
"10111010110101011101000101010111",
"11001110111011001110000010000000",
"10100110100110001001011111000011",
"00110110000011010011000110111001",
"10110100000101100011100101011101",
"10110011110111010000010010111101",
"00101000100000011011001001001101",
"00100011000111010101000000101111",
"11010101100000110001101010001110",
"10111001001000010010000010110011",
"00010000100001010010010111011011",
"11100101001110000111000100000010",
"10110110001111111101101111111000",
"00110000001111000100100001110111",
"01111010011001101100010010100001",
"01101011001010011011100110111001",
"10011100101101100110000111100000",
"01101111100010010010101110111001",
"11001100110000110111001100001110",
"10111000011000110010100100101001",
"11001000101000000000011101110111",
"01000001100011100000000001011001",
"01111100011111010000110000110100",
"10001001001000100100011100010111",
"11000110001000000110011111111110",
"11111110111100001011000000001000",
"10011000111000000111101011000000",
"01011000010100110000110101101111",
"11101110011000111001010101001110",
"00010011111001011010111111110010",
"11000010110011000011000011111001",
"11111001000111100010000011110100",
"10001001001110011011000101110101",
"01000010111001010110011011011011",
"10000011101000000111011000010110",
"11010101011010011001000000000011",
"00011001100100100110010110111110",
"11000100111100101011101110111100",
"10101001100010011111100000011100",
"00101111000000101101000110111000",
"11001110011110110111111010010110",
"00010111111101001110010110011101",
"10100110111100001001011000111001",
"11100000100101001110110100010100",
"01011100110111100101110110100100",
"11111110000000010101110000010001",
"01100110000000001010010010111011",
"01001010101100011011110100101001",
"01110001001100101010000111100111",
"01100110101000010000010100100101",
"00001111010010000001000100100111",
"00110110011110111010110110011110",
"11100100101100011010000100101011",
"11010001111110010100111111100011",
"01110111001011001111110100110001",
"01111011100000110100011111111111",
"00010110100100100110110110001010",
"01010010100101100010111001111000",
"00101110100001110101001100100111",
"10100001001001011101101000100101",
"10010000001011110101011111010001",
"10010110100001110110111100110101",
"11001111111101011000011001000101",
"00100111000000011110010001110110",
"00101101010111001101100111110101",
"10010101010011011100001101001011",
"10000011001100011000001100000100",
"10100100100101011101010001110011",
"00101011110100001101110000011111",
"10010000111101000111101011100100",
"11111101110010100010110000000010",
"00001000110101111010110110001010",
"11000111001010100101010000000010",
"00011111011010100001101100010100",
"00110111101001001010111010100110",
"00010111100101101001100100001111",
"11011000110010101000100011001011",
"10010100001010011010100011101110",
"00101101100001100011100111110100",
"11011000010111110010000110001011",
"11001001001110111110011111111011",
"01100010001000111100011110110011",
"01110101110000101100011010011011",
"10000011110010011100111001100100",
"10111010000110011000101011111000",
"01010011101111110101010010101001",
"10011110001011101111111111101011",
"10110010100000101100101011010000",
"00110011011111001100001100110110",
"10101100001010011111011011000110",
"10100000001001111101000010000110",
"11010111111110101101001011100101",
"00010011010110010110100000010001",
"10101011110101010000001010111010",
"11001011111010101000111001110011",
"00010010010111101010110110000010",
"10011110110011000000011010000001",
"00100110100010000101011001110000",
"11100110100110100100110101100011",
"11001101101001000101101001101100",
"00101111110101100011010101011110",
"00110110010101110111010011101111",
"00100110101101000100100010101010",
"10111010001000010100001101010011",
"10111111111011011001010001001110",
"00111010100101011010100011000000",
"01011110000111001001010000111001",
"01010010100110110001011101011001",
"01110001001111011011100000001101",
"11111110110001010000111000011111",
"10100100000101101101010001010110",
"01100011011010000011001101110000",
"10110111011100000011110001100111",
"01001011000001011111110001100001",
"11000010111110110111100001110000",
"11011001100000010011001001011111",
"00000110101101011101001000100011",
"10100000101101111000010101010100",
"01011001010100001110100101111100",
"01011000110001010111000010001111",
"01110010101000010001111110000111",
"11111100110111000100010011100101",
"00110010111000110000110100100010",
"11110000010000110101110001100100",
"01010110111100100000101101100101",
"00010111001010100101010111111111",
"00101110101000010000110011100000",
"10101111111100110111011110011100",
"01011000010101101101001000110001",
"11001000110011000100110111100011",
"10100011110001100010101111100101",
"11001100110011000011000101001011",
"00110001000111100001000100100011",
"11100110010111111100111101011011",
"00110011011000110010101101010011",
"11011010010001101001101010111110",
"10111010000110001111110101110111",
"10101011001111011011011001110000",
"00100101111000101100000001010000",
"10000100000000110010011011111111",
"01000000101101011110011001011011",
"10000101001110100110000100101100",
"01110011100110001111001101111101",
"00011010010101011011011100110000",
"01001110011111110110000000010011",
"11110101101100000110111110111110",
"10111101000110011100000001111110",
"01110011010100111110111011100110",
"11010100010001000001011001111110",
"01010111001000100011001100000011",
"11101011111110000111101010011101",
"10101111011110010000010100110101",
"01001010111100001110100101101000",
"10111010111010100101011111101101",
"11000101100000100010101100000101",
"01011010010000010011100000011111",
"11100000010001000111110111110000",
"00011000110110101010010100110000",
"00111111100011010110111010100100",
"00011000111100011001011011110101",
"01111100101001110010111100100010",
"00101010000001000110110110100111",
"01100111001011001111011111010011",
"01010111101010010000000001011100",
"10001000101100010100100001110010",
"10100000111010100001001000100110",
"00011010110100000100100000100100",
"11111100101010110000001010011011",
"11011000000010110010001001001111",
"01010110111011000011101010111010",
"00101011100000001111000011101000",
"01000010111011011111011101010100",
"00101111110111000010111011110000",
"10011100010010010101100001101000",
"10001100101011010010110011100100",
"11000110010011011100011000001111",
"01110100000010101110001101000110",
"11111010110111110100011011100110",
"00000000110000101111101000111001",
"11010010100100010111011101101110",
"10010011110111011001010101100001",
"01111000100111011110011000110000",
"00110101010101010001101011000011",
"01101110100000110111000100001000",
"01100000110101100000101110101011",
"00110110010100110001011011010100",
"01010111101100000111111010110100",
"10000010001100010100100101011010",
"01011001111111111011110110011110",
"10011100101100010001101101100001",
"11110110010010010001011000000110",
"00111101111011001110110001111001",
"11110100101110100001101000001101",
"00110001111101111100111110111111",
"01011011111111110111101000010001",
"01001110011101110100111000011001",
"00101110100100001111000101111111",
"01111100000111110100111101101011",
"01101011001101000110010111101010",
"00001000010011011111010011110110",
"01010110010011000011010010010010",
"00011111001001000100100101111111",
"00001100100111110100101101100110",
"01101100001011111000010001001110",
"00111001010110100110110110111100",
"00011101111110110101111100011101",
"11110101101100100000000110010101",
"11010100001011101100100110110000",
"10110011100111101110111000001110",
"10010000111000011010010101011110",
"00000101000011000001010111100100",
"01010001000001011110001101110101",
"00100011011110000100110001010011",
"00110101000000011101110001000100",
"01110110011100010010011010000110",
"10100101001011000111101110110011",
"11011100001000100111101001101000",
"01100110001100011110111000001100",
"00010010110110101100110101110001",
"00111001100110000001001110000000",
"01010110110101100110111011101111",
"00001110100111110111000101001100",
"00100110000001011000110111001101",
"00100111101110011100011001111101",
"01011001111100011001010001101001",
"01000010001011110100111110001111",
"00101110110110000010100001110011",
"00110101110110001010011010000010",
"00100101001101101110111010111001",
"11011001010100001111001011010101",
"01010101010100101011100100101001",
"11101111001010111111111001010100",
"11111010011111110011010011011100",
"10000010101111100101001000000001",
"00111101101111011011101011111011",
"11111100110000001011101110111111",
"10110110011001000101000011111000",
"01110011101010111110010000101011",
"01001001001111110001111001101001",
"00111100000011001110100111001010",
"01000101110100100110011001010110",
"11001010101011000101101100010110",
"00101011101111011111011101010010",
"10110110111111111100101110000101",
"11000010100101100001100001110001",
"00011101111111011001111010010101",
"10100001000101001011001100100010",
"01110111111011110011001011111110",
"00100100011101010100110110100100",
"01011100111001010011010001011001",
"01011010010011011111010000100110",
"10101110111101111011101110110101",
"11001001110001110100110110010100",
"10000100010010100111010011011110",
"01101111100110111000100110110111",
"10110100011101100000001101010111",
"10001000010001101000011000101000",
"11110010110100010110111110101001",
"00111011101000100110101000011110",
"00101110110111100101100101110011",
"10011001010000111110011001110111",
"10001000101010100010011001001110",
"11000101000000011101110111001001",
"10000110100000101000110101001111",
"00001100000001000111010010011111",
"10100100100000000010101111100100",
"01001111011101101011000101101001",
"10110100011101110000011000000000",
"00011111110010100101010110111001",
"11101001110111000010000110101111",
"11001010001011011111110001001010",
"11011001011101111010101101100110",
"10000101001110011101101010000110",
"00011111001100111100111001000110",
"01010111000111000000111110110110",
"10010111101000000000001100101100",
"10101111010000110001011110000010",
"00100110001111010100011001010000",
"00100010100000110110110001011010",
"00001001010000100101011000101110",
"10101001000001011111100110101001",
"11111011011000110000001101010011",
"01100100111011011001110000111100",
"01001010110110011011010010111100",
"11100100101111101110111101111110",
"11110000001000100101111111001110",
"01010101100100011000100110000010",
"10101101001011000011111011000100",
"11000011010000111101100000100100",
"10010100000100100101101110110001",
"10111100010011110001111000100011",
"00010000111011001101001010111110",
"00000100001101110001000101101001",
"11111011011110010011101110110111",
"11000000001100100011101010100011",
"10011101111111001010100000010001",
"11001010100010101110000101000000",
"00101001000010010001000011101000",
"01000101111011011110010010010011",
"00001000100010101001011000101000",
"00001111000000001100100011000000",
"10101011101010101000101001111101",
"01011100100011001111010000010110",
"11001000101110111100110010101110",
"01101011011001010111010101000001",
"01010001101001111001100000110111",
"01111101100101100011011111101100",
"10001101111101101011011001011011",
"11101111100001001000100111000011",
"00111101111111110111010110010101",
"01100110110000100011101101010011",
"00110101001101110011110110100000",
"01011100100010110000011100101010",
"10110000101100000111100101010111",
"01010111111101101100110000111110",
"11001001001010100010000101100101",
"10100010100000011010110101111110",
"00101011001000010010000001001001",
"10001110001000110011110011101110",
"00110011101010111011011001110001",
"00101010001110001000101001101100",
"00011110011101111000111111110100",
"00101000101101101101011000100100",
"11001000110001000111100001111011",
"10110010000011000101001000000000",
"00100101010100010110110010010001",
"00011100000001110011100110100111",
"00000001110111010011111011010101",
"01101101101011101101000111011110",
"11001010010001110100001001011100",
"11111000100010000001001001110101",
"00111001110010111100110000100000",
"11111010110101001110111100011110",
"11110101001010011000001101100110",
"10110000000011000010110010111110",
"10011101110100011100101110110101",
"00001110011001011100000000100011",
"11110101110010001001011111110011",
"00100000111101001111100010100100",
"11010111001111111111001110100111",
"01001100000101100001100011101101",
"11000101000110011000101010100001",
"11010001101101000000110001011011",
"11000010101101010111101101100001",
"10000100100001110101011010111001",
"00000111101111111110001100010101",
"01001101110001011101100111000001",
"10001000111011000111110010001010",
"10010111001101101100010011111110",
"00000011110000010110101110101000",
"01100111011011100100101001011101",
"00101011101101000000101001000110",
"11010100100110111111101000101000",
"11000011111101000000010111111000",
"01011001000101001010111000010001",
"00001101111111011100110111100001",
"11000001001010101110110111101100",
"10001111101010010111011010011001",
"10111010011001000111011110000101",
"11111110011000010010000110111101",
"01111001010010001110101100101000",
"10001101011101111110111010100101",
"01000111001100011001001000111101",
"10010101001010111111100110100001",
"10001000010111001000000000101001",
"01011100010001111000011100011111",
"10100101001010111101110000000010",
"01011001000110100110001111001010",
"00100100111000110011011011111111",
"00111110100010010000011110100111",
"11010110010110110011000111111011",
"00101000110011011101000100011001",
"10111111101100000011101000001111",
"00100111001011101111001011010111",
"11111101001011000001100101011110",
"11100100111010110011100011111101",
"01111010111101001011101001100110",
"11000000110110010000100001000001",
"11111100010011110111100111100100",
"01000111010101101100001001010000",
"11011110001001100001000101010000",
"11100110000010110101000010000110",
"11010111100100010011010011111001",
"01011001001011011010100101101100",
"11110001010001010000000111001011",
"10100000010111110011101110101001",
"00110001001001101100100100111110",
"10010010000100010111000000101011",
"10001101011011100101000001011101",
"11101100101001111110010111101110",
"00111010100111000100110001111000",
"11010011111001111110101110001111",
"01100111011101111011000110101101",
"11111011111000000110010100111110",
"11100100101000111100101100001011",
"11000111100010111000010100010111",
"01101100101100101000100011001100",
"01011110010010010010111111000101",
"10111110011011001101110000000110",
"11011101001110100010010011110011",
"10010111100110101000010101110011",
"01000110110010111010010011110111",
"10011110111101011101011011001010",
"11110111111100100110111000110110",
"10011011011000100110100010000010",
"01010011110101100110100001000100",
"10001000000010100100111001110001",
"11010111011111111111110110010000",
"00100000000010100100110100100000",
"00010011010101011011000001101001",
"11111010001000011011001010110001",
"11001110000001101111100100011010",
"01000001101011010011011111001001",
"01011001101011100001111101010010",
"01011011111010111010001000111000",
"11011001110100010011110111000111",
"11100011100011101110001101001001",
"01111101111010011001010000010100",
"00100001111110111011111101001111",
"01111011010100001110011011001011",
"01011101110011010110111001100110",
"11000010000111001000101111000010",
"00001000110110000101101010101001",
"10001011100001000100110101011100",
"00100100001110101100001100101100",
"11010010010001011000001011001110",
"10110111000100000001011110011110",
"00101001110001011000000001011110",
"10101011010110010010101101000111",
"10010101101001111000101100110011",
"01010111001101110010101000000011",
"11000111010101100011011101000100",
"11011111000110010100010010101001",
"01000001011101111110100111110101",
"01010100011110100111110111110010",
"01010110011100101001010001110001",
"00101110001010001001110101000100",
"00111010000110000101011011001000",
"00101000110010001010110100010010",
"10011101101001110011101000010001",
"11100111000000111111101110101011",
"01000101001011000110111000111001",
"11100010010101001110001001110110",
"10101110000010010001101011100101",
"01010000111001000000011100011101",
"10110110111000010111010110001110",
"01101010110010010100010000000010",
"11100010001100010100000100110001",
"10111101000011101100011011010000",
"00011101111100000010000010111101",
"10011011100001011110110010100101",
"01001001010010010100110000000100",
"01001101001110111100011101010011",
"01010111000100111010011101000010",
"10100111101010111111110100011111",
"10100110011001011111000100101100",
"00001110100110100111101101110100",
"00001101011010011110110011010111",
"01100000110001101011101001100110",
"00101110101101011001011110000010",
"10001110110011111101010101001011",
"11111110001011110110111010110101",
"01001101100011100110110010101111",
"01110101011010101001010100111111",
"00100000000011111010000001001001",
"01010110000000111001110000111110",
"01110011000010110111111101001110",
"00111001001101011000011010101111",
"01101100110001011101010011001100",
"11011111100110110111011111011011",
"01011010001000000001110111011101",
"11111010010000100111101000010111",
"00111010111001101101100001000011",
"01100101000000001110010000110001",
"01100000011010000111001111001101",
"11100011101001010001011101000000",
"00110000001101010111101111111100",
"11010100011010100001001011001010",
"10011111000110111110000000100111",
"01001000100110100111100010110011",
"10101000001111000001110010101011",
"11001110000100100101000110101010",
"10110111110100011110111101100000",
"01000110011011111111101011111010",
"11110001000001110111011000001111",
"00101111011000111011110101011010",
"11100000111100010000001111000010",
"10001001100000111101101100110111",
"10111011111000000000000100000110",
"00000101111001101100000010101110",
"11001101101111101101010101101101",
"11000010011010101011110011100011",
"01010000101011101111101111100100",
"11000001011101101111110011000001",
"00110001011110111101110101001011",
"10110011011100101111111101010010",
"10011101010011101001111000001101",
"00110111001111011001011101000001",
"10010101000110010000010011000011",
"11010100110001101111000010110011",
"00010110001010000010001000011111",
"10101011100000101010100001111010",
"10101100011111010110111111111110",
"00111100100110101110001111110001",
"10101001100110010101011100001000",
"11011101000111101010110001010000",
"11000101101110000101000111111110",
"01100011011001000111110101010111",
"11001000100110100110100101101110",
"11000101001101011101110000110011",
"01001110010110110110001010111000",
"01111100011100110111001101110101",
"00000101111001010000010000001001",
"01000010110110011100101000011110",
"00011100000011010010011000101000",
"10100110010011100100001101000101",
"10000010111000110111001110010110",
"00100001010011111101010111111000",
"00111100011010010000111110111110",
"00011110001111010011011010000111",
"01111001000000111111001110101111",
"00001001010001101001100110011010",
"01000010110011001011101101001011",
"10111001101101110010101100100111",
"01100011000111010111100110011000",
"11011101011000010101100011101110",
"11011011001000000101111111011111",
"00001101110000101000110010000110",
"10101001011100111100000101011111",
"11010011011110101101111010000100",
"01101001011100110111000000011010",
"11111101011011101000111100010010",
"10101110101010010100110001001110",
"11110110010100001001111100110101",
"01100101100010011111011101001001",
"11111100001101011010001100111110",
"00010000100101101110110100011011",
"11001101010101100010101111000011",
"10110110111001010011000001100001",
"11110000000101110100111000110011",
"01100111100001110111010110001100",
"10101100100000000101110111110001",
"00011011100011001010111110000000",
"10001000100011010001011011000000",
"01111101100000001101000111011001",
"10110100001001001001101000010100",
"11110010001001011010011111101111",
"11000001111001110010011010011010",
"01000001110101011110010101000001",
"11000100010000010010001000011110",
"00101011010010010101010101011011",
"11000111001110011011110101111000",
"10110011000100100001001110110001",
"00111101100010100101110010101101",
"10110011011101011001110001111101",
"10110001100001001011111101000110",
"01000100000011001000100110011001",
"00000001011001101000010101010111",
"00000101111111010001100110100101",
"10010011100011000110010011100011",
"11101010011000110001110111010110",
"00111110011110010001101110100100",
"00011110100001111011011111101010",
"01110010010011000001111111100001",
"01010001010110000110111011101010",
"00110100001000100000010100100010",
"11111010100011101010011001011111",
"11101111001101001001000001001001",
"11000001110010000110001111010111",
"10100111010010000011000010110010",
"00101001100111001011010000011110",
"01011010101111011100110100101111",
"00111110011011010101110110010011",
"01011001101011111111110001010101",
"00111111110100111110001011101011",
"00001011000101011000100111000010",
"00001011011101111000101000110000",
"11100110000010111101110110110111",
"10010010110100100110101100001111",
"00111001011001011110110010111100",
"01111101001101011000100011100101",
"10000001100000101111111001000110",
"10111111001110011100011110101000",
"10011001010001010011001110100111",
"11000000101110100111100111101101",
"00011010100011111010010101110011",
"01110100001001011111011010111100",
"00101100100010010110100001100010",
"01100001001100100010100101101101",
"00011001011011000011100101110111",
"10111111100111010101100011010100",
"10011001100100010011000100110101",
"01010010011011111100001111100100",
"11000110010000010111101011110011",
"11011001001101010011010111010110",
"11000111110001000111100100111001",
"00000011101101011101001100100010",
"10001100000010111000101110111111",
"00101011100110111011001001011101",
"01000111100101001101010110101011",
"00110011101101010000101000100010",
"00110000101001010100001010100101",
"11111001101000010011110000000000",
"11101010110100000010101101001011",
"00100110001010101010010001100010",
"11011010000011001011010100101100",
"11000000101110111001010101010010",
"00011001101010100000111000000000",
"01000101011110101101001100110000",
"00011111101001101001110111110101",
"00001011101111000100111000100011",
"00111000000111110100111011010010",
"00000100011010100101110100000100",
"00111011110101010010000111110100",
"00100111001000011010110001000111",
"00100011100001101001100111001000",
"10001110101100000101100100110011",
"11110010100110010001100101100101",
"01000001110100101110110110011100",
"11011101011110100101000111010100",
"10110010011000100011110100100011",
"01010000010111010011100000000101",
"11111001111101110001001011001110",
"11000001111000001101000011111111",
"01111100010110001111101000101010",
"00111011100000100000110011111111",
"10011101100110001101001001011001",
"10011001100110110100010100100111",
"00010111110011101011001111001000",
"11100000010100101000010001000011",
"10111000101010011111101001000101",
"10011000011100011101001100010110",
"00111001001010001000011000011000",
"10010010000111110011000100110010",
"11100000010010100011001001011111",
"10000110001000000010100000000011",
"00100110111111001111111000101011",
"01111000101110010100000101101000",
"10100010111100001101111111110000",
"11011100001011100100111101011111",
"01010101010100110001110100010011",
"10110010010000111000000101000111",
"11001000001000010011100111000010",
"01110100001001000101001001000111",
"00010011001000110010010101111110",
"01000111110100010111000011101000",
"00110000101110111111011111010111",
"11001001010011100001010000101001",
"10111010100101110101000000111100",
"10011011101000011111010011000001",
"00110010100101101001111111100011",
"10001110101111101001010100011111",
"10010010111010010010010000100110",
"00110111000110100111110001001101",
"10001010100011001011000011110010",
"11110000010000110000001001100110",
"11001110000001110111001110111101",
"01111110110011100101110011011100",
"01010100001001111001101111000000",
"10000111110001111011100000110110",
"10011100100000101100001010101110",
"00101010101110001001100000100110",
"00010110101111100101010100000001",
"00000010000010010011111000110111",
"11001001000000011101011001001000",
"10000010010111100000011111010100",
"00001011111000010011011110010110",
"00010101100000010010110101010010",
"01001001001111000110101001110000",
"00011111001111100010010111111011",
"10010010100010100111111010011001",
"01111110000111111001100001111110",
"11010001001011001010111001000001",
"00110000101101100011100001100001",
"10101000010011111011100101101010",
"10011001100100111101101110010001",
"01011111011010100011010110110111",
"10111000100110001100011001011010",
"11011000100010111100010101011101",
"10000110101000000011101000010111",
"11101110100111000100000000001011",
"00110101110000111001011011110111",
"01001101000110110010101100111011",
"11110000011111100010101010111101",
"11111110000110100000111011001100",
"10111001101110101001010100101101",
"01101001011101010000100011101010",
"11100011101100101001011101000011",
"01100111100101001010000101101000",
"10010111011110000010001000111110",
"10111111100100000001000000111110",
"10111111110001111101101110101000",
"01011100000011101010001100000101",
"11011100010111101011011000111000",
"10010100101001110110100101011111",
"01001010111001001000101000010101",
"10100000000101010111010000100101",
"10111001100000001100101000100000",
"10001111000110011011011001100000",
"00001001000110101010100100011010",
"01101110110110111110001110011100",
"00011101101110000010110001001110",
"01001101000111100011000110100110",
"11100010101001111100001100100111",
"00100001100001110011111101110010",
"11000100101100010100001011111011",
"00001010111111000100100001011100",
"11000001000001100101000100110100",
"10001100100001000101110111100110",
"01011000011111100111001101110011",
"11100011000110001111001100111010",
"11111100000110000000011001001110",
"10111111001001111001011000111111",
"01100110110001011111100111011111",
"11100110100000011001101000110010",
"00110001101010101000001111110100",
"00100110010101111010100111111001",
"00011000100011111010011000001001",
"10110101011100010110000001011001",
"11100101001001100001110001100010",
"01011011000111001001111100111101",
"00000010110111100100100010110000",
"01101100000100010110001100111110",
"00101111011111000111101010101111",
"01011110001110101111101110101000",
"10101110100010000110100000101011",
"11001101010001110100001110001110",
"11010000000011111010011110011101",
"00111001000100001110011011010001",
"11001001101000101001111110011100",
"00101001000001010111011001110111",
"11011000011110001001110101001101",
"11000010000000011001110011000101",
"10111111001111101001011100101101",
"10100010010101000101101100001111",
"00100010000111100001100011111100",
"01001000101011000000010100001000",
"00101011000100101010111101101010",
"00110100010001010010000101111010",
"10010000001110001100101111001100",
"01110111001001000111100110101011",
"11000111111011010111010011000101",
"01100011001101011101110011101001",
"10101100000101000101001100100101",
"11001111110100101011110110001111",
"01011010100111001011101101010001",
"00011111010011101100000000110100",
"00111010011111010010100011001111",
"01011000010111111010011100000101",
"11011111100110001010111010000011",
"11111000100001010110001110100001",
"10100101100001010011000111000000",
"01010011010101010010110010100111",
"10111001010111011101001101000000",
"10110010001111001110000000100111",
"11110010101100111100000101000100",
"01100101100001001001111101010010",
"10011101110001100111000010101110",
"00111000000010011110010101111001",
"10010110010101011100100001011011",
"00101111001011100101111100100101",
"00011011011100001111001111101001",
"00001011001001000001111101010110",
"01000111100001010100011100001110",
"10111111100000001111110111010111",
"11000111100001100100111101011100",
"01011110110011111011111000001011",
"11010110001010001010110000000000",
"11110101100010001110000001001011",
"00110101110000010101101010000100",
"01010010100001101011100000110110",
"01001000110010111000000100000110",
"00100101110110111110010011011110",
"10101110101100101100111010011111",
"10010101000110011001011010011101",
"10111110100110110101001110110111",
"01100000100010001110100101101011",
"11011111101001100010010000110011",
"11010011001111001010101010110000",
"00011000101010111000110000111000",
"10101100011111001101101010110100",
"11010000101101010111000110110010",
"11100100110001110110001110011111",
"01110110000011010101000111111101",
"10000000001110000101011110001000",
"01100000000110001010100011001111",
"10100000110110111101101100001111",
"00011111100110011010011010100110",
"01100110000111010010000110000101",
"01000110001111001001111010100100",
"10111100010001011100110110000110",
"00110110101011100000011001000100",
"10110011100001100111011010001000",
"00001001001101001011111001111010",
"00111111001111110000110111011111",
"00001001000001101110001111101000",
"11010111101001111101001000110110",
"00111101011100000110001000100000",
"11010101100111011001010101100110",
"11010110000110111110111001011001",
"10001001001001100111110100100001",
"00011111110010101101000110001010",
"01101101111011011110000011000000",
"00111010111010011111000000011110",
"01101001010110010110000010101101",
"00011011000000101001100011101101",
"00111000111111010011110111000111",
"00010100100000010011000010100110",
"10101101110111010111101111101000",
"00011010101101010000100100101011",
"10001001000111001010000010001010",
"11001100111000011001010000110111",
"01100101110000011110110010101111",
"11110011001010101110000101001100",
"11101110111010000110100111010000",
"00110000010001111101100101011000",
"11011111101101010110111110010010",
"10100000101000111101000110001011",
"01111001110101100100011000111110",
"11011011000010010001111000011101",
"10001100000110000011101101101101",
"01100101011100100110110000100010",
"10110010000100000010100001111010",
"11100000001111111111110111100001",
"10011011110010000011001010100100",
"00111100100101100010010001010010",
"01001100000100000000101111111101",
"10101110100100011001011110011101",
"10111011001000111101100000110011",
"10011111000101011010101100011010",
"11110110111110110011010100011010",
"01010110100100101101110111001110",
"11111000000111010010000000001101",
"00110101001011101000101001010110",
"11101101110101100100000101100010",
"10100110100100011011110010011000",
"01100110010100000011110000111000",
"11001101011011010001011100000111",
"01001011110000101010100001011010",
"00101001000001011000110100011001",
"00110101010010110001100110000001",
"10100011100000111001111001001010",
"11010111111111100001011011111011",
"00111100000000101010001011011110",
"00010101101111111100010110100011",
"01111110111010101011011000011111",
"01010101001011111101001100010101",
"11110101111001011110101100111001",
"10110100100011100110001011100111",
"01101010111111111100001010011010",
"00110010110101010011110010110111",
"00001110100111110001101000001111",
"00000010000001001000011001101010",
"11000011110011011010010001100101",
"00010101110101011000101001101001",
"10011010001010111000100011110111",
"01111100001001011100011010100001",
"10000010011010000011010110011100",
"10111111000101100101111010111001",
"10101011011011011100001010110101",
"01101101100111110111111001101110",
"11011001100101000010000101011010",
"11000101100111011001010101101001",
"00001010111110100010111010010100",
"10010001000110100000000010010100",
"11110010001010000101110010011011",
"00100101101000010000000100001000",
"11011000010100111100010111010110",
"00100100100010111011011100100111",
"11110000010100100101111110110101",
"11010101011001011010000011110011",
"00100100111000001100001010011100",
"10111010001010100000000000011010",
"10011111100101010100000101010010",
"01001000110010010001101000101001",
"00001110011100111111011011010100",
"00010111101111111010010110111011",
"10000001100111101111011011111110",
"11110000111001100110110001101001",
"00110011000011110001010100111010",
"10000011010010011110010010110111",
"01111001110110101010000000010101",
"10111101101011000110101100000011",
"11101010001011001111111111001010",
"00110010101011101010110011010011",
"11011101011011000001010101001011",
"01101100110110001010110011101101",
"01001010011110100101101010101011",
"01110111110100111110010110011101");

  signal op1,op2,ans1,ans,answ,low,high: std_logic_vector(31 downto 0);
  signal addr: std_logic_vector(19 downto 0) := (others=>'0');
  signal miss: std_logic_vector(31 downto 0) := (others=>'0');
  signal rom_o: std_logic_vector(7 downto 0) := (others=>'1');
  signal uart_go: std_logic;
  signal uart_busy: std_logic := '0';
  signal iter: std_logic_vector(31 downto 0) := (others=>'0');
  signal state: std_logic_vector(4 downto 0) := (others=>'0');
  signal state2: std_logic_vector(4 downto 0) := (others=>'0');

begin

  ib: IBUFG port map (
   i=>MCLK1,
   o=>iclk);
  bg: BUFG port map (
    i=>iclk,
    o=>clk);

  fmuler:fmul port map
    (clk, op1, op2, ans);

  rs232c: u232c generic map (wtime=>x"1ADB")
  port map (
    clk=>clk,
    data=>rom_o,
    go=>uart_go,
    busy=>uart_busy,
    tx=>rs_tx);


 cal: process(clk)
 begin
   if rising_edge(clk) then-- hoge clk後に返答
     if state = "00000" then
       state<=state+1;
       addr<=addr+3;
       op1<=rom(conv_integer(addr));
       op2<=rom(conv_integer(addr+1));
       ans1<=rom(conv_integer(addr+2));
     elsif state = "00001" then
       state<=state+1;
     elsif state = "00010" then
       state<=state+1;
       answ<=ans;
       state2<="00000";
     elsif state = "00011" and uart_go = '1'then --op1の出力
       state2<=state2+1;
       if op1(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "00100" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "00101" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "00110" and uart_go = '1'then --op2の出力
       state2<=state2+1;
       if op2(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "00111" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01000" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01001" and uart_go = '1'then --outputの出力
       state2<=state2+1;
       if answ(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01010" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01011" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01100" and uart_go = '1'then --answerの出力
       state2<=state2+1;
       if ans1(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01101" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01110" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01111" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10000" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10001" then --low,highとの比較
       state<=state+1;
       low<=ans1 - 3;
     elsif state = "10010" then
       state<=state+1;
       high<=ans1 + 3;
     elsif state = "10011" then
       iter<=iter+1;
       state<=state+1;
       if high < answ or low > answ then
         miss<=miss+1;
       end if;
     elsif state = "10100" and uart_go = '1'then --iterの出力
       state2<=state2+1;
       if iter(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "10101" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10110" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10111" and uart_go = '1'then --missの出力
       state2<=state2+1;
       if miss(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "11000" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11001" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "11010" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11011" and uart_go = '1'then
       state<="00000";
       rom_o<=x"0a";
     end if;
   end if;
 end process;

    send_msg: process(clk)
  begin
    if rising_edge(clk) then
      if uart_busy='0' and uart_go='0' then
        uart_go<='1';
      else
        uart_go<='0';
      end if;
    end if;
  end process;
  
end VHDL;
