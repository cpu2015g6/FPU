/home/mizuta1018/HW/FPU/VHDL/fsin/fsin.vhd