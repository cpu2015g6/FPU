/home/mizuta1018/HW/FPU/VHDL/fsin/fmul_2.vhd