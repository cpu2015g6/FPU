/home/mizuta1018/HW/FPU/VHDL/fmul/octmul.vhd