/home/mizuta1018/HW/FPU/VHDL/fadd/u232c.vhd