/home/mizuta1018/HW/FPU/VHDL/fsin/fadd_2.vhd