/home/mizuta1018/HW/FPU/VHDL/finv/finv.vhd