library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity blockram is

  generic (
    dwidth : integer := 13;
    awidth : integer := 10);

  port (
    clk  : in  std_logic;
    we   : in  std_logic;
    di   : in  std_logic_vector(dwidth - 1 downto 0);
    do   : out std_logic_vector(dwidth - 1 downto 0);
    addr : in  std_logic_vector(awidth - 1 downto 0));

end entity;

architecture behavioral of blockram is

  type ram_type is
    array(0 to (2 ** awidth) - 1) of std_logic_vector(dwidth - 1 downto 0);

  signal ram : ram_type := ("0110101000001",
"0110100110101",
"0110100101010",
"0110100011111",
"0110100010100",
"0110100001001",
"0110011111101",
"0110011110010",
"0110011100111",
"0110011011100",
"0110011010001",
"0110011000110",
"0110010111011",
"0110010110000",
"0110010100110",
"0110010011011",
"0110010010000",
"0110010000101",
"0110001111010",
"0110001110000",
"0110001100101",
"0110001011010",
"0110001010000",
"0110001000101",
"0110000111010",
"0110000110000",
"0110000100101",
"0110000011011",
"0110000010000",
"0110000000110",
"0101111111100",
"0101111110001",
"0101111100111",
"0101111011101",
"0101111010010",
"0101111001000",
"0101110111110",
"0101110110100",
"0101110101001",
"0101110011111",
"0101110010101",
"0101110001011",
"0101110000001",
"0101101110111",
"0101101101101",
"0101101100011",
"0101101011001",
"0101101001111",
"0101101000101",
"0101100111011",
"0101100110001",
"0101100101000",
"0101100011110",
"0101100010100",
"0101100001010",
"0101100000001",
"0101011110111",
"0101011101101",
"0101011100100",
"0101011011010",
"0101011010000",
"0101011000111",
"0101010111101",
"0101010110100",
"0101010101010",
"0101010100001",
"0101010010111",
"0101010001110",
"0101010000100",
"0101001111011",
"0101001110010",
"0101001101000",
"0101001011111",
"0101001010110",
"0101001001101",
"0101001000011",
"0101000111010",
"0101000110001",
"0101000101000",
"0101000011111",
"0101000010110",
"0101000001100",
"0101000000011",
"0100111111010",
"0100111110001",
"0100111101000",
"0100111011111",
"0100111010110",
"0100111001101",
"0100111000101",
"0100110111100",
"0100110110011",
"0100110101010",
"0100110100001",
"0100110011000",
"0100110010000",
"0100110000111",
"0100101111110",
"0100101110101",
"0100101101101",
"0100101100100",
"0100101011011",
"0100101010011",
"0100101001010",
"0100101000010",
"0100100111001",
"0100100110000",
"0100100101000",
"0100100011111",
"0100100010111",
"0100100001111",
"0100100000110",
"0100011111110",
"0100011110101",
"0100011101101",
"0100011100101",
"0100011011100",
"0100011010100",
"0100011001100",
"0100011000011",
"0100010111011",
"0100010110011",
"0100010101011",
"0100010100010",
"0100010011010",
"0100010010010",
"0100010001010",
"0100010000010",
"0100001111010",
"0100001110010",
"0100001101001",
"0100001100001",
"0100001011001",
"0100001010001",
"0100001001001",
"0100001000001",
"0100000111001",
"0100000110010",
"0100000101010",
"0100000100010",
"0100000011010",
"0100000010010",
"0100000001010",
"0100000000010",
"0011111111011",
"0011111110011",
"0011111101011",
"0011111100011",
"0011111011011",
"0011111010100",
"0011111001100",
"0011111000100",
"0011110111101",
"0011110110101",
"0011110101101",
"0011110100110",
"0011110011110",
"0011110010111",
"0011110001111",
"0011110000111",
"0011110000000",
"0011101111000",
"0011101110001",
"0011101101001",
"0011101100010",
"0011101011011",
"0011101010011",
"0011101001100",
"0011101000100",
"0011100111101",
"0011100110110",
"0011100101110",
"0011100100111",
"0011100100000",
"0011100011000",
"0011100010001",
"0011100001010",
"0011100000010",
"0011011111011",
"0011011110100",
"0011011101101",
"0011011100110",
"0011011011110",
"0011011010111",
"0011011010000",
"0011011001001",
"0011011000010",
"0011010111011",
"0011010110100",
"0011010101101",
"0011010100101",
"0011010011110",
"0011010010111",
"0011010010000",
"0011010001001",
"0011010000010",
"0011001111011",
"0011001110101",
"0011001101110",
"0011001100111",
"0011001100000",
"0011001011001",
"0011001010010",
"0011001001011",
"0011001000100",
"0011000111101",
"0011000110111",
"0011000110000",
"0011000101001",
"0011000100010",
"0011000011011",
"0011000010101",
"0011000001110",
"0011000000111",
"0011000000001",
"0010111111010",
"0010111110011",
"0010111101101",
"0010111100110",
"0010111011111",
"0010111011001",
"0010111010010",
"0010111001011",
"0010111000101",
"0010110111110",
"0010110111000",
"0010110110001",
"0010110101011",
"0010110100100",
"0010110011110",
"0010110010111",
"0010110010001",
"0010110001010",
"0010110000100",
"0010101111101",
"0010101110111",
"0010101110000",
"0010101101010",
"0010101100100",
"0010101011101",
"0010101010111",
"0010101010001",
"0010101001010",
"0010101000100",
"0010100111110",
"0010100110111",
"0010100110001",
"0010100101011",
"0010100100100",
"0010100011110",
"0010100011000",
"0010100010010",
"0010100001100",
"0010100000101",
"0010011111111",
"0010011111001",
"0010011110011",
"0010011101101",
"0010011100111",
"0010011100000",
"0010011011010",
"0010011010100",
"0010011001110",
"0010011001000",
"0010011000010",
"0010010111100",
"0010010110110",
"0010010110000",
"0010010101010",
"0010010100100",
"0010010011110",
"0010010011000",
"0010010010010",
"0010010001100",
"0010010000110",
"0010010000000",
"0010001111010",
"0010001110100",
"0010001101110",
"0010001101000",
"0010001100010",
"0010001011101",
"0010001010111",
"0010001010001",
"0010001001011",
"0010001000101",
"0010000111111",
"0010000111001",
"0010000110100",
"0010000101110",
"0010000101000",
"0010000100010",
"0010000011101",
"0010000010111",
"0010000010001",
"0010000001011",
"0010000000110",
"0010000000000",
"0001111111010",
"0001111110101",
"0001111101111",
"0001111101001",
"0001111100100",
"0001111011110",
"0001111011000",
"0001111010011",
"0001111001101",
"0001111001000",
"0001111000010",
"0001110111100",
"0001110110111",
"0001110110001",
"0001110101100",
"0001110100110",
"0001110100001",
"0001110011011",
"0001110010110",
"0001110010000",
"0001110001011",
"0001110000101",
"0001110000000",
"0001101111010",
"0001101110101",
"0001101101111",
"0001101101010",
"0001101100101",
"0001101011111",
"0001101011010",
"0001101010100",
"0001101001111",
"0001101001010",
"0001101000100",
"0001100111111",
"0001100111010",
"0001100110100",
"0001100101111",
"0001100101010",
"0001100100100",
"0001100011111",
"0001100011010",
"0001100010100",
"0001100001111",
"0001100001010",
"0001100000101",
"0001011111111",
"0001011111010",
"0001011110101",
"0001011110000",
"0001011101011",
"0001011100101",
"0001011100000",
"0001011011011",
"0001011010110",
"0001011010001",
"0001011001100",
"0001011000110",
"0001011000001",
"0001010111100",
"0001010110111",
"0001010110010",
"0001010101101",
"0001010101000",
"0001010100011",
"0001010011110",
"0001010011001",
"0001010010011",
"0001010001110",
"0001010001001",
"0001010000100",
"0001001111111",
"0001001111010",
"0001001110101",
"0001001110000",
"0001001101011",
"0001001100110",
"0001001100001",
"0001001011100",
"0001001011000",
"0001001010011",
"0001001001110",
"0001001001001",
"0001001000100",
"0001000111111",
"0001000111010",
"0001000110101",
"0001000110000",
"0001000101011",
"0001000100110",
"0001000100010",
"0001000011101",
"0001000011000",
"0001000010011",
"0001000001110",
"0001000001001",
"0001000000101",
"0001000000000",
"0000111111011",
"0000111110110",
"0000111110001",
"0000111101101",
"0000111101000",
"0000111100011",
"0000111011110",
"0000111011010",
"0000111010101",
"0000111010000",
"0000111001100",
"0000111000111",
"0000111000010",
"0000110111101",
"0000110111001",
"0000110110100",
"0000110101111",
"0000110101011",
"0000110100110",
"0000110100001",
"0000110011101",
"0000110011000",
"0000110010100",
"0000110001111",
"0000110001010",
"0000110000110",
"0000110000001",
"0000101111101",
"0000101111000",
"0000101110011",
"0000101101111",
"0000101101010",
"0000101100110",
"0000101100001",
"0000101011101",
"0000101011000",
"0000101010100",
"0000101001111",
"0000101001011",
"0000101000110",
"0000101000010",
"0000100111101",
"0000100111001",
"0000100110100",
"0000100110000",
"0000100101011",
"0000100100111",
"0000100100010",
"0000100011110",
"0000100011001",
"0000100010101",
"0000100010001",
"0000100001100",
"0000100001000",
"0000100000011",
"0000011111111",
"0000011111011",
"0000011110110",
"0000011110010",
"0000011101101",
"0000011101001",
"0000011100101",
"0000011100000",
"0000011011100",
"0000011011000",
"0000011010011",
"0000011001111",
"0000011001011",
"0000011000111",
"0000011000010",
"0000010111110",
"0000010111010",
"0000010110101",
"0000010110001",
"0000010101101",
"0000010101001",
"0000010100100",
"0000010100000",
"0000010011100",
"0000010011000",
"0000010010011",
"0000010001111",
"0000010001011",
"0000010000111",
"0000010000011",
"0000001111110",
"0000001111010",
"0000001110110",
"0000001110010",
"0000001101110",
"0000001101010",
"0000001100101",
"0000001100001",
"0000001011101",
"0000001011001",
"0000001010101",
"0000001010001",
"0000001001101",
"0000001001000",
"0000001000100",
"0000001000000",
"0000000111100",
"0000000111000",
"0000000110100",
"0000000110000",
"0000000101100",
"0000000101000",
"0000000100100",
"0000000100000",
"0000000011100",
"0000000011000",
"0000000010100",
"0000000010000",
"0000000001100",
"0000000001000",
"0000000000100",
"0000000000000",
"1111111110000",
"1111111100000",
"1111111010000",
"1111111000000",
"1111110110000",
"1111110100000",
"1111110010001",
"1111110000001",
"1111101110001",
"1111101100010",
"1111101010010",
"1111101000011",
"1111100110011",
"1111100100100",
"1111100010101",
"1111100000101",
"1111011110110",
"1111011100111",
"1111011011000",
"1111011001001",
"1111010111001",
"1111010101010",
"1111010011011",
"1111010001100",
"1111001111110",
"1111001101111",
"1111001100000",
"1111001010001",
"1111001000010",
"1111000110100",
"1111000100101",
"1111000010110",
"1111000001000",
"1110111111001",
"1110111101011",
"1110111011100",
"1110111001110",
"1110110111111",
"1110110110001",
"1110110100011",
"1110110010100",
"1110110000110",
"1110101111000",
"1110101101010",
"1110101011100",
"1110101001110",
"1110101000000",
"1110100110010",
"1110100100100",
"1110100010110",
"1110100001000",
"1110011111010",
"1110011101100",
"1110011011110",
"1110011010001",
"1110011000011",
"1110010110101",
"1110010101000",
"1110010011010",
"1110010001100",
"1110001111111",
"1110001110001",
"1110001100100",
"1110001010110",
"1110001001001",
"1110000111100",
"1110000101110",
"1110000100001",
"1110000010100",
"1110000000111",
"1101111111001",
"1101111101100",
"1101111011111",
"1101111010010",
"1101111000101",
"1101110111000",
"1101110101011",
"1101110011110",
"1101110010001",
"1101110000100",
"1101101110111",
"1101101101011",
"1101101011110",
"1101101010001",
"1101101000100",
"1101100111000",
"1101100101011",
"1101100011110",
"1101100010010",
"1101100000101",
"1101011111001",
"1101011101100",
"1101011100000",
"1101011010011",
"1101011000111",
"1101010111010",
"1101010101110",
"1101010100010",
"1101010010110",
"1101010001001",
"1101001111101",
"1101001110001",
"1101001100101",
"1101001011001",
"1101001001100",
"1101001000000",
"1101000110100",
"1101000101000",
"1101000011100",
"1101000010000",
"1101000000100",
"1100111111000",
"1100111101101",
"1100111100001",
"1100111010101",
"1100111001001",
"1100110111101",
"1100110110010",
"1100110100110",
"1100110011010",
"1100110001111",
"1100110000011",
"1100101110111",
"1100101101100",
"1100101100000",
"1100101010101",
"1100101001001",
"1100100111110",
"1100100110010",
"1100100100111",
"1100100011100",
"1100100010000",
"1100100000101",
"1100011111010",
"1100011101110",
"1100011100011",
"1100011011000",
"1100011001101",
"1100011000001",
"1100010110110",
"1100010101011",
"1100010100000",
"1100010010101",
"1100010001010",
"1100001111111",
"1100001110100",
"1100001101001",
"1100001011110",
"1100001010011",
"1100001001000",
"1100000111101",
"1100000110011",
"1100000101000",
"1100000011101",
"1100000010010",
"1100000000111",
"1011111111101",
"1011111110010",
"1011111100111",
"1011111011101",
"1011111010010",
"1011111000111",
"1011110111101",
"1011110110010",
"1011110101000",
"1011110011101",
"1011110010011",
"1011110001000",
"1011101111110",
"1011101110011",
"1011101101001",
"1011101011111",
"1011101010100",
"1011101001010",
"1011101000000",
"1011100110101",
"1011100101011",
"1011100100001",
"1011100010111",
"1011100001100",
"1011100000010",
"1011011111000",
"1011011101110",
"1011011100100",
"1011011011010",
"1011011010000",
"1011011000110",
"1011010111100",
"1011010110010",
"1011010101000",
"1011010011110",
"1011010010100",
"1011010001010",
"1011010000000",
"1011001110110",
"1011001101100",
"1011001100010",
"1011001011001",
"1011001001111",
"1011001000101",
"1011000111011",
"1011000110010",
"1011000101000",
"1011000011110",
"1011000010101",
"1011000001011",
"1011000000001",
"1010111111000",
"1010111101110",
"1010111100101",
"1010111011011",
"1010111010001",
"1010111001000",
"1010110111110",
"1010110110101",
"1010110101100",
"1010110100010",
"1010110011001",
"1010110001111",
"1010110000110",
"1010101111101",
"1010101110011",
"1010101101010",
"1010101100001",
"1010101010111",
"1010101001110",
"1010101000101",
"1010100111100",
"1010100110011",
"1010100101001",
"1010100100000",
"1010100010111",
"1010100001110",
"1010100000101",
"1010011111100",
"1010011110011",
"1010011101010",
"1010011100001",
"1010011011000",
"1010011001111",
"1010011000110",
"1010010111101",
"1010010110100",
"1010010101011",
"1010010100010",
"1010010011001",
"1010010010000",
"1010010000111",
"1010001111110",
"1010001110110",
"1010001101101",
"1010001100100",
"1010001011011",
"1010001010010",
"1010001001010",
"1010001000001",
"1010000111000",
"1010000110000",
"1010000100111",
"1010000011110",
"1010000010110",
"1010000001101",
"1010000000100",
"1001111111100",
"1001111110011",
"1001111101011",
"1001111100010",
"1001111011010",
"1001111010001",
"1001111001001",
"1001111000000",
"1001110111000",
"1001110101111",
"1001110100111",
"1001110011111",
"1001110010110",
"1001110001110",
"1001110000101",
"1001101111101",
"1001101110101",
"1001101101100",
"1001101100100",
"1001101011100",
"1001101010100",
"1001101001011",
"1001101000011",
"1001100111011",
"1001100110011",
"1001100101011",
"1001100100010",
"1001100011010",
"1001100010010",
"1001100001010",
"1001100000010",
"1001011111010",
"1001011110010",
"1001011101010",
"1001011100010",
"1001011011010",
"1001011010001",
"1001011001001",
"1001011000001",
"1001010111010",
"1001010110010",
"1001010101010",
"1001010100010",
"1001010011010",
"1001010010010",
"1001010001010",
"1001010000010",
"1001001111010",
"1001001110010",
"1001001101011",
"1001001100011",
"1001001011011",
"1001001010011",
"1001001001011",
"1001001000100",
"1001000111100",
"1001000110100",
"1001000101100",
"1001000100101",
"1001000011101",
"1001000010101",
"1001000001110",
"1001000000110",
"1000111111110",
"1000111110111",
"1000111101111",
"1000111101000",
"1000111100000",
"1000111011000",
"1000111010001",
"1000111001001",
"1000111000010",
"1000110111010",
"1000110110011",
"1000110101011",
"1000110100100",
"1000110011100",
"1000110010101",
"1000110001110",
"1000110000110",
"1000101111111",
"1000101110111",
"1000101110000",
"1000101101001",
"1000101100001",
"1000101011010",
"1000101010011",
"1000101001011",
"1000101000100",
"1000100111101",
"1000100110101",
"1000100101110",
"1000100100111",
"1000100100000",
"1000100011000",
"1000100010001",
"1000100001010",
"1000100000011",
"1000011111100",
"1000011110100",
"1000011101101",
"1000011100110",
"1000011011111",
"1000011011000",
"1000011010001",
"1000011001010",
"1000011000011",
"1000010111011",
"1000010110100",
"1000010101101",
"1000010100110",
"1000010011111",
"1000010011000",
"1000010010001",
"1000010001010",
"1000010000011",
"1000001111100",
"1000001110101",
"1000001101110",
"1000001101000",
"1000001100001",
"1000001011010",
"1000001010011",
"1000001001100",
"1000001000101",
"1000000111110",
"1000000110111",
"1000000110001",
"1000000101010",
"1000000100011",
"1000000011100",
"1000000010101",
"1000000001111",
"1000000001000",
"1000000000001",
"0111111111010",
"0111111110100",
"0111111101101",
"0111111100110",
"0111111011111",
"0111111011001",
"0111111010010",
"0111111001011",
"0111111000101",
"0111110111110",
"0111110110111",
"0111110110001",
"0111110101010",
"0111110100100",
"0111110011101",
"0111110010110",
"0111110010000",
"0111110001001",
"0111110000011",
"0111101111100",
"0111101110110",
"0111101101111",
"0111101101001",
"0111101100010",
"0111101011100",
"0111101010101",
"0111101001111",
"0111101001000",
"0111101000010",
"0111100111011",
"0111100110101",
"0111100101110",
"0111100101000",
"0111100100010",
"0111100011011",
"0111100010101",
"0111100001111",
"0111100001000",
"0111100000010",
"0111011111011",
"0111011110101",
"0111011101111",
"0111011101001",
"0111011100010",
"0111011011100",
"0111011010110",
"0111011001111",
"0111011001001",
"0111011000011",
"0111010111101",
"0111010110110",
"0111010110000",
"0111010101010",
"0111010100100",
"0111010011110",
"0111010010111",
"0111010010001",
"0111010001011",
"0111010000101",
"0111001111111",
"0111001111001",
"0111001110011",
"0111001101100",
"0111001100110",
"0111001100000",
"0111001011010",
"0111001010100",
"0111001001110",
"0111001001000",
"0111001000010",
"0111000111100",
"0111000110110",
"0111000110000",
"0111000101010",
"0111000100100",
"0111000011110",
"0111000011000",
"0111000010010",
"0111000001100",
"0111000000110",
"0111000000000",
"0110111111010",
"0110111110100",
"0110111101110",
"0110111101000",
"0110111100010",
"0110111011101",
"0110111010111",
"0110111010001",
"0110111001011",
"0110111000101",
"0110110111111",
"0110110111001",
"0110110110100",
"0110110101110",
"0110110101000",
"0110110100010",
"0110110011100",
"0110110010111",
"0110110010001",
"0110110001011",
"0110110000101",
"0110101111111",
"0110101111010",
"0110101110100",
"0110101101110",
"0110101101001",
"0110101100011",
"0110101011101",
"0110101010111",
"0110101010010",
"0110101001100",
"0110101000110");

  signal reg_addr : std_logic_vector(awidth - 1 downto 0);

begin

  process(clk)
  begin
    if rising_edge(clk) then
      if we = '1' then
        ram(conv_integer(addr)) <= di;
      end if;
      reg_addr <= addr;
    end if;
  end process;

  do <= ram(conv_integer(reg_addr));

end behavioral;
