library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity invblockram2 is

  generic (
    dwidth : integer := 13;
    awidth : integer := 10);

  port (
    clk  : in  std_logic;
    we   : in  std_logic;
    di   : in  std_logic_vector(dwidth - 1 downto 0);
    do   : out std_logic_vector(dwidth - 1 downto 0);
    addr : in  std_logic_vector(awidth - 1 downto 0));

end invblockram2;

architecture behavioral of invblockram2 is

  type ram_type is
    array(0 to (2 ** awidth) - 1) of std_logic_vector(dwidth - 1 downto 0);

  signal ram : ram_type := ("1111111110011",
"1111111010000",
"1111110110000",
"1111110010010",
"1111101110011",
"1111101010011",
"1111100110001",
"1111100010011",
"1111011110100",
"1111011010101",
"1111010110101",
"1111010011000",
"1111001111001",
"1111001011010",
"1111000111001",
"1111000011100",
"1110111111101",
"1110111011111",
"1110111000000",
"1110110100000",
"1110110000100",
"1110101100101",
"1110101001000",
"1110100101010",
"1110100001011",
"1110011101101",
"1110011001111",
"1110010110010",
"1110010010100",
"1110001111001",
"1110001011011",
"1110000111101",
"1110000100000",
"1110000000000",
"1101111100110",
"1101111001010",
"1101110101010",
"1101110010000",
"1101101110010",
"1101101010110",
"1101100111000",
"1101100011101",
"1101100000000",
"1101011100100",
"1101011001001",
"1101010101011",
"1101010010000",
"1101001110100",
"1101001011001",
"1101000111011",
"1101000100000",
"1101000000110",
"1100111101010",
"1100111001110",
"1100110110010",
"1100110010110",
"1100101111101",
"1100101100000",
"1100101000100",
"1100100101010",
"1100100001111",
"1100011110101",
"1100011011001",
"1100010111110",
"1100010100100",
"1100010001010",
"1100001101111",
"1100001010101",
"1100000111010",
"1100000100000",
"1100000000101",
"1011111101100",
"1011111010010",
"1011110110111",
"1011110011110",
"1011110000100",
"1011101101001",
"1011101010000",
"1011100110110",
"1011100011100",
"1011100000100",
"1011011101001",
"1011011010000",
"1011010110111",
"1011010100000",
"1011010000101",
"1011001101011",
"1011001010011",
"1011000111010",
"1011000100000",
"1011000000110",
"1010111101111",
"1010111010110",
"1010110111101",
"1010110100110",
"1010110001101",
"1010101110011",
"1010101011011",
"1010101000100",
"1010100101010",
"1010100010011",
"1010011111010",
"1010011100010",
"1010011001001",
"1010010110011",
"1010010011011",
"1010010000000",
"1010001101011",
"1010001010010",
"1010000111100",
"1010000100100",
"1010000001110",
"1001111110110",
"1001111011110",
"1001111000111",
"1001110101111",
"1001110010111",
"1001110000000",
"1001101101010",
"1001101010011",
"1001100111100",
"1001100100110",
"1001100001110",
"1001011110110",
"1001011100000",
"1001011001011",
"1001010110011",
"1001010011110",
"1001010000110",
"1001001101111",
"1001001011010",
"1001001000011",
"1001000101101",
"1001000011000",
"1001000000000",
"1000111101010",
"1000111010101",
"1000110111111",
"1000110101001",
"1000110010100",
"1000110000000",
"1000101101000",
"1000101010010",
"1000100111011",
"1000100100101",
"1000100010010",
"1000011111011",
"1000011100110",
"1000011010010",
"1000010111011",
"1000010100110",
"1000010010000",
"1000001111101",
"1000001100110",
"1000001010010",
"1000000111101",
"1000000101000",
"1000000010100",
"1000000000000",
"0111111101001",
"0111111010101",
"0111111000000",
"0111110101010",
"0111110011000",
"0111110000000",
"0111101101111",
"0111101011010",
"0111101000110",
"0111100110000",
"0111100011101",
"0111100001010",
"0111011110100",
"0111011100000",
"0111011001100",
"0111010111000",
"0111010100100",
"0111010010001",
"0111001111101",
"0111001101000",
"0111001010110",
"0111001000000",
"0111000101101",
"0111000011010",
"0111000000111",
"0110111110010",
"0110111100000",
"0110111001101",
"0110110111010",
"0110110100101",
"0110110010011",
"0110110000000",
"0110101101100",
"0110101011001",
"0110101000101",
"0110100110010",
"0110100100000",
"0110100001100",
"0110011111011",
"0110011101000",
"0110011010101",
"0110011000011",
"0110010101111",
"0110010011100",
"0110010001010",
"0110001111001",
"0110001100100",
"0110001010011",
"0110001000000",
"0110000101110",
"0110000011100",
"0110000001010",
"0101111110111",
"0101111100101",
"0101111010010",
"0101111000000",
"0101110101110",
"0101110011100",
"0101110001011",
"0101101111001",
"0101101100111",
"0101101010110",
"0101101000100",
"0101100110001",
"0101100011111",
"0101100001101",
"0101011111101",
"0101011101011",
"0101011011001",
"0101011001001",
"0101010110101",
"0101010100011",
"0101010010100",
"0101010000000",
"0101001110000",
"0101001100000",
"0101001001111",
"0101000111101",
"0101000101011",
"0101000011011",
"0101000001010",
"0100111111001",
"0100111100110",
"0100111010110",
"0100111000110",
"0100110110101",
"0100110100100",
"0100110010100",
"0100110000000",
"0100101110011",
"0100101100000",
"0100101010000",
"0100101000000",
"0100100110000",
"0100100011111",
"0100100001111",
"0100100000000",
"0100011101110",
"0100011011110",
"0100011001101",
"0100010111011",
"0100010101101",
"0100010011100",
"0100010001011",
"0100010000000",
"0100001101100",
"0100001011011",
"0100001001100",
"0100000111011",
"0100000101101",
"0100000011100",
"0100000001110",
"0100000000000",
"0011111101100",
"0011111011101",
"0011111001101",
"0011110111101",
"0011110101110",
"0011110011101",
"0011110001110",
"0011110000000",
"0011101110000",
"0011101100000",
"0011101010000",
"0011101000000",
"0011100110001",
"0011100100011",
"0011100010100",
"0011100000110",
"0011011110100",
"0011011100110",
"0011011010110",
"0011011001000",
"0011010111001",
"0011010101010",
"0011010011001",
"0011010001011",
"0011010000000",
"0011001101101",
"0011001011110",
"0011001010000",
"0011001000000",
"0011000110010",
"0011000100011",
"0011000010101",
"0011000001000",
"0010111111000",
"0010111101000",
"0010111011001",
"0010111001101",
"0010110111101",
"0010110101111",
"0010110100000",
"0010110010010",
"0010110000101",
"0010101110101",
"0010101100110",
"0010101010111",
"0010101001100",
"0010100111100",
"0010100101110",
"0010100100000",
"0010100010010",
"0010100000110",
"0010011110110",
"0010011101000",
"0010011011001",
"0010011001100",
"0010010111110",
"0010010101111",
"0010010100010",
"0010010010100",
"0010010001000",
"0010001111000",
"0010001101011",
"0010001011100",
"0010001010000",
"0010001000000",
"0010000110011",
"0010000100101",
"0010000011001",
"0010000001011",
"0010000000000",
"0001111110000",
"0001111100010",
"0001111010110",
"0001111001001",
"0001110111011",
"0001110101101",
"0001110100000",
"0001110010100",
"0001110000110",
"0001101111001",
"0001101101010",
"0001101011101",
"0001101010001",
"0001101000011",
"0001100110111",
"0001100101001",
"0001100011101",
"0001100010000",
"0001100000100",
"0001011110110",
"0001011101000",
"0001011011100",
"0001011010000",
"0001011000100",
"0001010110100",
"0001010101000",
"0001010011100",
"0001010001111",
"0001010000000",
"0001001110110",
"0001001101001",
"0001001011100",
"0001001010001",
"0001001000100",
"0001000110110",
"0001000101011",
"0001000011101",
"0001000010000",
"0001000000101",
"0000111111000",
"0000111101101",
"0000111100000",
"0000111010011",
"0000111001000",
"0000110111100",
"0000110101110",
"0000110100011",
"0000110011000",
"0000110001011",
"0000110000000",
"0000101110010",
"0000101100110",
"0000101011011",
"0000101001111",
"0000101000011",
"0000100110111",
"0000100101010",
"0000100011101",
"0000100010011",
"0000100000111",
"0000011111010",
"0000011101111",
"0000011100010",
"0000011011000",
"0000011001100",
"0000011000000",
"0000010110101",
"0000010101001",
"0000010011101",
"0000010010001",
"0000010000101",
"0000001111010",
"0000001101110",
"0000001100011",
"0000001011000",
"0000001001101",
"0000001000000",
"0000000110100",
"0000000101010",
"0000000011101",
"0000000010011",
"0000000001000",
"0000000000000",
"1111111100010",
"1111111001100",
"1111110110010",
"1111110100000",
"1111110001010",
"1111101110010",
"1111101011010",
"1111101000110",
"1111100101110",
"1111100011000",
"1111100000000",
"1111011101110",
"1111011011000",
"1111011000000",
"1111010101100",
"1111010010110",
"1111001111110",
"1111001100110",
"1111001010100",
"1111001000000",
"1111000101000",
"1111000010010",
"1111000000000",
"1110111101000",
"1110111010000",
"1110110111100",
"1110110100110",
"1110110010000",
"1110101111010",
"1110101100110",
"1110101010010",
"1110100111010",
"1110100101000",
"1110100010100",
"1110100000000",
"1110011101000",
"1110011010010",
"1110010111110",
"1110010101010",
"1110010010010",
"1110001111110",
"1110001101010",
"1110001010100",
"1110001000000",
"1110000101100",
"1110000010110",
"1110000000000",
"1101111110000",
"1101111011100",
"1101111001000",
"1101110110010",
"1101110011010",
"1101110001000",
"1101101110100",
"1101101100000",
"1101101001110",
"1101100110110",
"1101100100100",
"1101100001110",
"1101100000000",
"1101011101010",
"1101011010100",
"1101011000000",
"1101010101100",
"1101010011000",
"1101010000000",
"1101001101110",
"1101001011100",
"1101001001000",
"1101000110110",
"1101000100000",
"1101000001110",
"1101000000000",
"1100111100100",
"1100111010010",
"1100111000000",
"1100110101100",
"1100110011010",
"1100110001000",
"1100101110010",
"1100101100000",
"1100101001110",
"1100100111000",
"1100100100110",
"1100100010100",
"1100100000000",
"1100011101110",
"1100011100011",
"1100011010000",
"1100010111101",
"1100010101010",
"1100010010111",
"1100010000101",
"1100001110010",
"1100001011111",
"1100001001101",
"1100000111010",
"1100000100111",
"1100000010101",
"1100000000010",
"1011111110000",
"1011111011101",
"1011111001011",
"1011110111000",
"1011110100110",
"1011110010100",
"1011110000001",
"1011101101111",
"1011101011101",
"1011101001011",
"1011100111001",
"1011100100110",
"1011100010100",
"1011100000010",
"1011011110000",
"1011011011110",
"1011011001100",
"1011010111010",
"1011010101001",
"1011010010111",
"1011010000101",
"1011001110011",
"1011001100001",
"1011001010000",
"1011000111110",
"1011000101100",
"1011000011011",
"1011000001001",
"1010111111000",
"1010111100110",
"1010111010101",
"1010111000011",
"1010110110010",
"1010110100000",
"1010110001111",
"1010101111110",
"1010101101101",
"1010101011011",
"1010101001010",
"1010100111001",
"1010100101000",
"1010100010111",
"1010100000110",
"1010011110101",
"1010011100011",
"1010011010011",
"1010011000010",
"1010010110001",
"1010010100000",
"1010010001111",
"1010001111110",
"1010001101101",
"1010001011101",
"1010001001100",
"1010000111011",
"1010000101010",
"1010000011010",
"1010000001001",
"1001111111001",
"1001111101000",
"1001111011000",
"1001111000111",
"1001110110111",
"1001110100110",
"1001110010110",
"1001110000101",
"1001101110101",
"1001101100101",
"1001101010101",
"1001101000100",
"1001100110100",
"1001100100100",
"1001100010100",
"1001100000100",
"1001011110100",
"1001011100100",
"1001011010011",
"1001011000011",
"1001010110100",
"1001010100100",
"1001010010100",
"1001010000100",
"1001001110100",
"1001001100100",
"1001001010100",
"1001001000101",
"1001000110101",
"1001000100101",
"1001000010101",
"1001000000110",
"1000111110110",
"1000111100111",
"1000111010111",
"1000111000111",
"1000110111000",
"1000110101000",
"1000110011001",
"1000110001010",
"1000101111010",
"1000101101011",
"1000101011011",
"1000101001100",
"1000100111101",
"1000100101110",
"1000100011110",
"1000100001111",
"1000100000000",
"1000011110001",
"1000011100010",
"1000011010011",
"1000011000100",
"1000010110101",
"1000010100110",
"1000010010111",
"1000010001000",
"1000001111001",
"1000001101010",
"1000001011011",
"1000001001100",
"1000000111101",
"1000000101110",
"1000000100000",
"1000000010001",
"1000000000010",
"0111111110100",
"0111111100101",
"0111111010110",
"0111111001000",
"0111110111001",
"0111110101010",
"0111110011100",
"0111110001101",
"0111101111111",
"0111101110001",
"0111101100010",
"0111101010100",
"0111101000101",
"0111100110111",
"0111100101001",
"0111100011010",
"0111100001100",
"0111011111110",
"0111011110000",
"0111011100001",
"0111011010011",
"0111011000101",
"0111010110111",
"0111010101001",
"0111010011011",
"0111010001101",
"0111001111111",
"0111001110001",
"0111001100011",
"0111001010101",
"0111001000111",
"0111000111001",
"0111000101011",
"0111000011101",
"0111000001111",
"0111000000010",
"0110111110100",
"0110111100110",
"0110111011000",
"0110111001011",
"0110110111101",
"0110110101111",
"0110110100010",
"0110110010100",
"0110110000110",
"0110101111001",
"0110101101011",
"0110101011110",
"0110101010000",
"0110101000011",
"0110100110101",
"0110100101000",
"0110100011011",
"0110100001101",
"0110100000000",
"0110011110011",
"0110011100101",
"0110011011000",
"0110011001011",
"0110010111101",
"0110010110000",
"0110010100011",
"0110010010110",
"0110010001001",
"0110001111100",
"0110001101110",
"0110001100001",
"0110001010100",
"0110001000111",
"0110000111010",
"0110000101101",
"0110000100000",
"0110000010011",
"0110000000110",
"0101111111010",
"0101111101101",
"0101111100000",
"0101111010011",
"0101111000110",
"0101110111001",
"0101110101101",
"0101110100000",
"0101110010011",
"0101110000110",
"0101101111010",
"0101101101101",
"0101101100000",
"0101101010100",
"0101101000111",
"0101100111011",
"0101100101110",
"0101100100010",
"0101100010101",
"0101100001001",
"0101011111100",
"0101011110000",
"0101011100011",
"0101011010111",
"0101011001011",
"0101010111110",
"0101010110010",
"0101010100101",
"0101010011001",
"0101010001101",
"0101010000001",
"0101001110100",
"0101001101000",
"0101001011100",
"0101001010000",
"0101001000100",
"0101000111000",
"0101000101011",
"0101000011111",
"0101000010011",
"0101000000111",
"0100111111011",
"0100111101111",
"0100111100011",
"0100111010111",
"0100111001011",
"0100110111111",
"0100110110011",
"0100110101000",
"0100110011100",
"0100110010000",
"0100110000100",
"0100101111000",
"0100101101100",
"0100101100001",
"0100101010101",
"0100101001001",
"0100100111101",
"0100100110010",
"0100100100110",
"0100100011010",
"0100100001111",
"0100100000011",
"0100011111000",
"0100011101100",
"0100011100000",
"0100011010101",
"0100011001001",
"0100010111110",
"0100010110010",
"0100010100111",
"0100010011011",
"0100010010000",
"0100010000101",
"0100001111001",
"0100001101110",
"0100001100010",
"0100001010111",
"0100001001100",
"0100001000001",
"0100000110101",
"0100000101010",
"0100000011111",
"0100000010100",
"0100000001000",
"0011111111101",
"0011111110010",
"0011111100111",
"0011111011100",
"0011111010001",
"0011111000101",
"0011110111010",
"0011110101111",
"0011110100100",
"0011110011001",
"0011110001110",
"0011110000011",
"0011101111000",
"0011101101101",
"0011101100010",
"0011101011000",
"0011101001101",
"0011101000010",
"0011100110111",
"0011100101100",
"0011100100001",
"0011100010110",
"0011100001100",
"0011100000001",
"0011011110110",
"0011011101011",
"0011011100001",
"0011011010110",
"0011011001011",
"0011011000001",
"0011010110110",
"0011010101011",
"0011010100001",
"0011010010110",
"0011010001011",
"0011010000001",
"0011001110110",
"0011001101100",
"0011001100001",
"0011001010111",
"0011001001100",
"0011001000010",
"0011000110111",
"0011000101101",
"0011000100011",
"0011000011000",
"0011000001110",
"0011000000011",
"0010111111001",
"0010111101111",
"0010111100100",
"0010111011010",
"0010111010000",
"0010111000110",
"0010110111011",
"0010110110001",
"0010110100111",
"0010110011101",
"0010110010010",
"0010110001000",
"0010101111110",
"0010101110100",
"0010101101010",
"0010101100000",
"0010101010110",
"0010101001100",
"0010101000010",
"0010100110111",
"0010100101101",
"0010100100011",
"0010100011001",
"0010100001111",
"0010100000101",
"0010011111100",
"0010011110010",
"0010011101000",
"0010011011110",
"0010011010100",
"0010011001010",
"0010011000000",
"0010010110110",
"0010010101101",
"0010010100011",
"0010010011001",
"0010010001111",
"0010010000101",
"0010001111100",
"0010001110010",
"0010001101000",
"0010001011110",
"0010001010101",
"0010001001011",
"0010001000001",
"0010000111000",
"0010000101110",
"0010000100101",
"0010000011011",
"0010000010001",
"0010000001000",
"0001111111110",
"0001111110101",
"0001111101011",
"0001111100010",
"0001111011000",
"0001111001111",
"0001111000101",
"0001110111100",
"0001110110010",
"0001110101001",
"0001110100000",
"0001110010110",
"0001110001101",
"0001110000011",
"0001101111010",
"0001101110001",
"0001101100111",
"0001101011110",
"0001101010101",
"0001101001100",
"0001101000010",
"0001100111001",
"0001100110000",
"0001100100111",
"0001100011101",
"0001100010100",
"0001100001011",
"0001100000010",
"0001011111001",
"0001011110000",
"0001011100111",
"0001011011101",
"0001011010100",
"0001011001011",
"0001011000010",
"0001010111001",
"0001010110000",
"0001010100111",
"0001010011110",
"0001010010101",
"0001010001100",
"0001010000011",
"0001001111010",
"0001001110001",
"0001001101000",
"0001001011111",
"0001001010110",
"0001001001110",
"0001001000101",
"0001000111100",
"0001000110011",
"0001000101010",
"0001000100001",
"0001000011001",
"0001000010000",
"0001000000111",
"0000111111110",
"0000111110101",
"0000111101101",
"0000111100100",
"0000111011011",
"0000111010011",
"0000111001010",
"0000111000001",
"0000110111001",
"0000110110000",
"0000110100111",
"0000110011111",
"0000110010110",
"0000110001101",
"0000110000101",
"0000101111100",
"0000101110100",
"0000101101011",
"0000101100011",
"0000101011010",
"0000101010010",
"0000101001001",
"0000101000001",
"0000100111000",
"0000100110000",
"0000100100111",
"0000100011111",
"0000100010110",
"0000100001110",
"0000100000110",
"0000011111101",
"0000011110101",
"0000011101101",
"0000011100100",
"0000011011100",
"0000011010100",
"0000011001011",
"0000011000011",
"0000010111011",
"0000010110010",
"0000010101010",
"0000010100010",
"0000010011010",
"0000010010001",
"0000010001001",
"0000010000001",
"0000001111001",
"0000001110001",
"0000001101000",
"0000001100000",
"0000001011000",
"0000001010000",
"0000001001000",
"0000001000000",
"0000000111000",
"0000000110000",
"0000000101000",
"0000000100000",
"0000000011000",
"0000000010000",
"0000000001000");

  signal reg_addr : std_logic_vector(awidth - 1 downto 0);

begin

  process(clk)
  begin
    if rising_edge(clk) then
      if we = '1' then
        ram(conv_integer(addr)) <= di;
      end if;
      reg_addr <= addr;
    end if;
  end process;

  do <= ram(conv_integer(reg_addr));

end behavioral;
