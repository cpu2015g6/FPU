/home/mizuta1018/HW/FPU/VHDL/fadd/revfadd.vhd