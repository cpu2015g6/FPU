/home/mizuta1018/HW/FPU/VHDL/fcos/absfadd.vhd