/home/mizuta1018/HW/FPU/VHDL/fsin/fmul_4.vhd