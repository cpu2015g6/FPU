library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity fputop is
  port(MCLK1: in std_logic;
       RS_TX: out std_logic);
  end fputop;

architecture VHDL of fputop is

component u232c
  generic (wtime: std_logic_vector(15 downto 0) := x"1ADB");
  Port ( clk  : in  STD_LOGIC;
         data : in  STD_LOGIC_VECTOR (7 downto 0);
         go   : in  STD_LOGIC;
         busy : out STD_LOGIC;
         tx   : out STD_LOGIC);
end component;

component finv
  port(clk: in std_logic;
		 op: in std_logic_vector(31 downto 0);
		 ans: out std_logic_vector(31 downto 0));
		 end component;

  signal clk,iclk: std_logic;
  type rom_t is array(0 to 3945) of std_logic_vector(31 downto 0);
  constant rom: rom_t := ("11100000000110000110011010111101",
"10011110110101110000001011100010",
"10110010010100100000101010100111",
"11001100100111000000000111010111",
"10001011111010001011111110011001",
"11110011000011001100100110000110",
"11011110101000111110010000111110",
"10100000010001111110111111100100",
"11011101010000000111000100110101",
"10100001101010100100011001000101",
"10111010100101100001101010110001",
"11000100010110100100110100110101",
"11001010010100001111101000101110",
"10110100100111001100110100111111",
"11101001001101110011100100011110",
"10010101101100101101011110010010",
"11010111011001000111000010001011",
"10100111100011110111000101010110",
"11000000101110010011111010101100",
"10111110001100001110001111100111",
"11010101001100000000111100111111",
"10101001101110100001111001101100",
"10110101010001100011000111000001",
"11001001101001010101010100101001",
"10011101110000000110010111111111",
"11100001001010100101000000110001",
"10101000111011101011101011110011",
"11010110000010010100001001101111",
"00011100110011011101000111100011",
"01100010000111110011010100001001",
"00111101101000100011001011001010",
"01000001010010100000011000110010",
"10101000101111001001000100011110",
"11010110001011011100011000011111",
"00000011110000000100101010011000",
"01111011001010100110100001110110",
"10111111011111001010010010101001",
"10111111100000011011001101100001",
"01011001010110101111101111000101",
"00100101100101011010001100001001",
"01111001000010110011111001110100",
"00000101111010110101001111110111",
"11000110010100000101010000011000",
"10111000100111010100101001000001",
"11001010111110100101100001110011",
"10110100000000101110010000100000",
"11011100111100110000101101000110",
"10100010000001101101001011000100",
"01001111101010101110010001001110",
"00101111001111111011111100111110",
"11011011101010001010110101110001",
"10100011010000100100001110100010",
"00001010010001110110000010011010",
"01110100101001000101101000000111",
"10010010110001110100011111000000",
"11101100001001000110111010000110",
"00010100000111111010010010001001",
"01101010110011010100001000100011",
"10010110010010010011111001111010",
"11101000101000101101001111000010",
"01000100101111010010010001100100",
"00111010001011010011111011010000",
"10011101011101100110001110101000",
"11100001100001001111111000101000",
"11110100110110100010101011011110",
"10001010000101100011001001010010",
"01100100110011100101100101011100",
"00011010000111101100110010000100",
"11010111000001011100011110101011",
"10100111111101001111000010000110",
"11110001111000010001110010011000",
"10001101000100011001000000110100",
"11000000000111000000111101100100",
"10111110110100011111100001101010",
"00111011000010101110000001100110",
"01000011111010111111001101010111",
"01001000100011110000110000101010",
"00110110011001010001001000011100",
"11001111001100100011010100110000",
"10101111101101111110000000010001",
"01011010011111000110110010100111",
"00100100100000011101000000101000",
"00110101001001101001100011001101",
"01001001110001001011000010111011",
"10000001100000010101110001100100",
"11111101011111010100111010001101",
"00101000111110011011011100011100",
"01010110000000110011100010110001",
"01111010001100111011001111000100",
"00000100101101100101100010011011",
"11101011101101100000110000100011",
"10010011001100111111111101000000",
"11011011001100001001000100000011",
"10100011101110011001010110100011",
"11111110000011101010010001001011",
"10000000111001011011100011101011",
"11100110000111110111100000011100",
"10011000110011010111101101010010",
"10011110001111111110001010000101",
"11100000101010101100010011100011",
"11000000101101101001010101111000",
"10111110001100110111011111011101",
"01011010011110110101101110001011",
"00100100100000100101110100110100",
"11001100111111000111010000101000",
"10110010000000011100110001001100",
"10011101111000011011111110000111",
"11100001000100010010011100100101",
"10100000001111000000000010100110",
"11011110101011100100101110100111",
"10111001110000110011100111101110",
"11000101001001111101100010100100",
"01000110100011011000101010000010",
"00111000011001111000001001000010",
"01100111111111000010000110110101",
"00010111000000011111011010111110",
"10111000001100000001000000010011",
"11000110101110100001110110001100",
"11011111110110011000000111000100",
"10011111000101101010011100010111",
"10101100101001001100101010010010",
"11010010010001101101100001110000",
"11010100101110111111110110110010",
"10101010001011100100111001100100",
"00101001111010000000000100110110",
"01010101000011010011110100001110",
"00001101100100000110110010000101",
"01110001011000101110001100111101",
"11111000000000001011010110010110",
"10000110111111101001011011010100",
"11011000010010001110001011011001",
"10100110101000110001111000000111",
"01001111000110011010011011011010",
"00101111110101010100001011101111",
"11101000000000100100110100010010",
"10010110111110110111101010101010",
"00111010110100001101011101010101",
"01000100000111001110011101101001",
"11011010000011110101101100011000",
"10100100111001001001001111111100",
"00000010111101101011101100000110",
"01111100000001001100111100010000",
"11100011011111011110001111111111",
"10011011100000010001000000111111",
"01101000101010111100110010000000",
"00010110001111101011110000010110",
"11111011111010001011010110001101",
"10000011000011001100111110011010",
"11001110000100011011011111101001",
"10110000111000001101111101000001",
"00010100000101001101110000101100",
"01101010110111000010000001010000",
"11010100011100101010111100110100",
"10101010100001110000010111101010",
"00100101011010011111000101011001",
"01011001100011000001000110000110",
"00100011101011000100111110101101",
"01011011001111100010101011100011",
"11000110100000101001010000100110",
"10111000011110101111000111000111",
"00000001010000010101111111011100",
"01111101101010010111010000100000",
"01101110001010010001011001100100",
"00010000110000011100101100001111",
"11000100000100001100111000000010",
"10111010111000100100101001111101",
"10111101010101100110110100010111",
"11000001100110001101000100110100",
"11011110011010011011000100101111",
"10100000100011000011011111111011",
"11110011011101011011011010011010",
"10001011100001010101101111010011",
"00111000000000101010110111001010",
"01000110111110101100000010001010",
"01001100010100110100100011110001",
"00110010100110110001011011010011",
"01110010101000011000111010101100",
"00001100010010101101001101101011",
"01101001001100111100100010001111",
"00010101101101100100001110000100",
"01000010110100010110100001011101",
"00111100000111000111101010111110",
"10111011011010011100100100010010",
"11000011100011000010100110100111",
"11100110000110010111111010011011",
"10011000110101010111101011011010",
"00010101100111101100011111111011",
"01101001010011100101111101000000",
"00010011110011100001100001001010",
"01101011000111101111111010100111",
"00100101011100101101001110001100",
"01011001100001101111000110110101",
"01111010111011001101001100100010",
"00000100000010100101110100101010",
"01100101011010100111111011011100",
"00011001100010111011110011111111",
"11101001110001110100110101100111",
"10010101001001000110100111011100",
"10111101110111110100011001111011",
"11000001000100101100001010110001",
"10111010001001101011010000100010",
"11000100110001001001000001111100",
"00101001100100010110101011001100",
"01010101011000010101011010000000",
"10001000010010001001011110101111",
"11110110101000110101101100100110",
"00010010110101111101110000110111",
"01101100000101111100110101001100",
"00111110001000001011001000111011",
"01000000110010111110100110100111",
"00111011100111010110110011110010",
"01000011010100000010011000101111",
"01111001010101000100100110000010",
"00000101100110100101101101100010",
"10011000001101100011001000101001",
"11100110101100111101100110101111",
"11010111110110101111000001101111",
"10100111000101011010101011001001",
"11101001001100111001011001100110",
"10010101101101100111011001101101",
"00001001111101100101011001000111",
"01110101000001010000010101100001",
"10000000101110001000000011011111",
"11111110001100011001100111011111",
"10100010010000100101001111100010",
"11011100101010001001111101010110",
"01000011111000001100101010001101",
"00111011000100011100010101010101",
"00001000111000111110101110101110",
"01110110000011111100010011110100",
"11010100001110101001111111100001",
"10101010101011111001010100011110",
"10110011000101010000111000011101",
"11001011110110111101011010001111",
"10110101001101000000000110111101",
"11001001101101100000100110011111",
"01110011101100001011111001101011",
"00001011001110010110010111110110",
"00110110010001111100110000101001",
"01001000101001000000000110001101",
"11000100000101111000001010111011",
"10111010110110000100011001110100",
"10110010110000111000101100111111",
"11001100001001111001001011010111",
"01101000111011000110111100011111",
"00010110000010101001011110110001",
"00011100110110011001010001011011",
"01100010000101101001101000111000",
"11111000110011101011011110001101",
"10000110000111101000010000101000",
"00101100011100000110100001001000",
"01010010100010000100110101001111",
"10010100101100111001010010110011",
"11101010001101100111100000100111",
"10000111101010000011011100111101",
"11110111010000101100110000100100",
"00010011010010111110100011100011",
"01101011101000001011001011010110",
"11000010111111111000100111011111",
"10111100000000000011101100101100",
"01001101010010010001001011010010",
"00110001101000101111011100011100",
"01011111001110100111010001100010",
"00011111101011111011111000010100",
"00010101000001100011010001101110",
"01101001111101000010101000000101",
"10111011101110111100011010111101",
"11000011001011101000000101101000",
"01011100011110100101010000010100",
"00100010100000101110011001101001",
"10111010100010000110001101111111",
"11000100011100000100000100101100",
"01100011111010001100110000000001",
"00011011000011001100001000000101",
"01011101111111011010001100001101",
"00100001000000010011000101001011",
"00111000010001011010110000100111",
"01000110101001011100010011101000",
"00001101100111001001101010101110",
"01110001010100010011110110101001",
"00000000111001000110001000101001",
"01111110000011110111101001011111",
"00110011110110010111000110001001",
"01001011000101101011001001010110",
"01100111001101011110110000011110",
"00010111101101000001111011101110",
"11001100100011011101111101110001",
"10110010011001101111011110101001",
"10000111000010101010101010010001",
"11110111111011000100111011110001",
"10010110101100011010100110010010",
"11101000001110000111000010010001",
"10100110110001111001001100010001",
"11011000001001000011000001111000",
"11010100101100011101111001010011",
"10101010001110000011100111011101",
"00001010010110101001010000010101",
"01110100100101011110101000000101",
"11000100100001001011101001011000",
"10111010011101101110000110001010",
"00000010011100010011011111110110",
"01111100100001111101011111110101",
"10000111011001101011111011111001",
"11110111100011100000001001001100",
"01101100010110010000110010010110",
"00010010100101101111100001101100",
"10110011001011110011111100010111",
"11001011101110101111101101111110",
"01100000001110111001100101101110",
"00011110101011101010101110001110",
"11010101101100110001110001110010",
"10101001001101101111001010101001",
"11111010110110001101110010111100",
"10000100000101110001100110111100",
"01110110101101111111001001110011",
"00001000001100100010001101100001",
"01000101000011100011011011000001",
"00111001111001100110100111011100",
"01011100100100001001110111011011",
"00100010011000101001010111010110",
"01010010110100110011101100110101",
"00101100000110110010000011101000",
"10100000011011001001111010110110",
"11011110100010100111101111010001",
"11101001001011100110010101100011",
"10010101101110111110010011101000",
"00110101011010001001010111000110",
"01001001100011001110001011010111",
"10000101100011000010001000011010",
"11111001011010011101010110101100",
"01011010010111011110000110100001",
"00100100100100111010111010111010",
"01111000111110100110110111110111",
"00000110000000101101100011100001",
"11101110010101110101111000001000",
"10010000100110000010011000111101",
"11000111001010010000001010100000",
"10110111110000011110000110111001",
"00001001111100100011001101001011",
"01110101000001110100101011111110",
"11100010010100100111011011100101",
"10011100100110111011000110011011",
"00001000100001001001011110100101",
"01110110011101110010001000100110",
"01101001001100011101110110111000",
"00010101101110000011101001111110",
"10111111001110100001110001111100",
"10111111101100000001000100010100",
"01000010100000100101101111111101",
"00111100011110110101110111100011",
"01111010010110001111010111001100",
"00000100100101110000100001001000",
"00001111000011010000000111000110",
"01101111111010000110001011000000",
"10001110111100000110010101111001",
"11110000000010000100111011100111",
"00001111111001000001000110001011",
"01101111000011111010110100010110",
"11101011110001000110000010100001",
"10010011001001101101110011000010",
"00111110010001100100101101011111",
"01000000101001010011111111001110",
"00011101011011011000110110110110",
"01100001100010011111000001111110",
"00100111111001101110001011011101",
"01010111000011011110110000111001",
"10011100100101000011001111100011",
"11100010010111010001101001000101",
"00101101010010111000100011011101",
"01010001101000001111111010100110",
"10010110011101001000000110001100",
"11101000100001100000010001100011",
"10000110001010111011011011101011",
"11111000101111101101010000001111",
"11101100110010010101001101100101",
"10010010001000101100001011010111",
"10011110001101011010001101001010",
"11100000101101000110011100100110",
"10011101100111011010100100011101",
"11100001010011111101011011000000",
"11000111110011100010101000111001",
"10110111000111101111000011010010",
"11110110000011011001011001111001",
"10001000111001110110111010110001",
"10110010101111000011001101101011",
"11001100001011100001110010100011",
"01001111000101101001001100101000",
"00101111110110011001111010001111",
"11001001010101101111011100110011",
"10110101100110000110111100000101",
"01011000000100000111100010011100",
"00100110111000101101000001000000",
"00000000111111010011011000001100",
"01111110000000010110100011101001",
"10111110110111011111101111101000",
"11000000000100111001110100111111",
"10000001010000101111001000010000",
"11111101101010000001011010000100",
"10010111111100111111111001100110",
"11100111000001100100110001101100",
"00000001111110001001011011111010",
"01111101000000111101000011001001",
"10111110001011000111101010110000",
"11000000101111011111101101110110",
"11001101011000011001100100100100",
"10110001100100010011111111011000",
"01110111100000011110001010001001",
"00000111011111000100100011101111",
"01010110111110010011110111110111",
"00101000000000110111100001111001",
"01001100010011110011101110110101",
"00110010100111100001111100010001",
"00101101000101100010101010001111",
"01010001110110100011011000100100",
"01110101101000101001010000110000",
"00001001010010011000110100101010",
"01000111010110101100111000100001",
"00110111100101011100001001000000",
"00100010011100101010001011110000",
"01011100100001110000110010111110",
"00011000010011110000011111100110",
"01100110100111100100011010100011",
"01110000000000010010000111011110",
"00001110111111011100000101011001",
"00101001011101010110101000010111",
"01010101100001011000010101100110",
"10110010100111110011001110011010",
"11001100010011011101001110111110",
"00011111110100101000111011011100",
"01011111000110111001111111100010",
"01101111110100011110100001110000",
"00001111000111000001101101000101",
"00111100101111000001100001111001",
"01000010001011100011010110010100",
"00001000111101001101011110100010",
"01110110000001011101010101000100",
"10101000110010101011111000000010",
"11010110001000011001111110111100",
"11001001010111011000011010101000",
"10110101100100111110101101100000",
"10110111011101101100101111100101",
"11000111100001001100010111111100",
"11010110010001100000111100110001",
"10101000101001010111001000000011",
"00111001000100010011100101010010",
"01000101111000011010001101000110",
"00001111100000110101111101011011",
"01101111011110010110110110011110",
"01110011001110111100110110101110",
"00001011101011100111101011110101",
"10111001001101101010010110100010",
"11000101101100110110011111111011",
"01010100100000010000001101111011",
"00101010011111011111110100011110",
"10100100000101010111100000110110",
"11011010110110110011101010000011",
"01100110001101100110100100111110",
"00011000101100111010001101100000",
"01010010010100101001101111100100",
"00101100100110111001011001000001",
"01010001000110101110001000111010",
"00101101110100111001000010110001",
"01010111001100000111110010111010",
"00100111101110011010101011111000",
"10111011001101011000100100011111",
"11000011101101001000000100101000",
"01101110111111111001100111110011",
"00010000000000000011001100011011",
"10010111000000011011010010011010",
"11100111111111001010001001000111",
"00101110010000110001100011100010",
"01010000101001111111010100010010",
"00100101010001111111111111100000",
"01011001101000111101011100100100",
"11100110000000000111010111101110",
"10011000111111110001010011111101",
"00011111111110011010011010101000",
"01011111000000110100000101010111",
"01011100100111011100011001111101",
"00100010010011111011000000001110",
"00111100011110010011001100101001",
"01000010100000110111111000101100",
"10111011110111000101110000000011",
"11000011000101001011001111011000",
"10001101001110111101000000111000",
"11110001101011100111100010011001",
"10000101010011011100100011111100",
"11111001100111110011101111101101",
"01110011110110010011010011100000",
"00001011000101101101110001101100",
"00010110011001001011101100101111",
"01101000100011110100001010000111",
"10110010111001111101100001100110",
"11001100000011010101010111101011",
"10111110110110011011011101010111",
"11000000000101101000001000000101",
"00001110001000110011101101001100",
"01110000110010001011111011010011",
"10101000000010000110100001101110",
"11010110111100000011100001111100",
"01010100010011111011011100100011",
"00101010100111011100000100011100",
"10010010011011001011001110110011",
"11101100100010100110111110001010",
"10111101100111111101001110000100",
"11000001010011010000010111001101",
"00101110011000110001011000111111",
"01010000100100000100110000010100",
"01010001101010010110110100111101",
"00101101010000010110011110111000",
"10110110110010011100011001110110",
"11001000001000100110011000000101",
"11100110100111100000111001001010",
"10011000010011110101000110110101",
"10011111000111001101011100001100",
"11011111110100001110110100011111",
"01010010100101111111011010110010",
"00101100010101111010000101101001",
"01100111010011000001011111111010",
"00010111101000001000110111000010",
"11111100000010110000010011101001",
"10000010111010111011010101011111",
"10001011011001010100001010101101",
"11110011100011101110110111011100",
"01101011010001100000101100010010",
"00010011101001010111010101110101",
"10011101000100000011111011010101",
"11100001111000110010101100011010",
"11111000000110000100101101001110",
"10000110110101110010100110011101",
"00011110100011100011011001000110",
"01100000011001100110101010100011",
"10011011011001000010100010010011",
"11100011100011111001111010010101",
"11000101111111111011100101110101",
"10111001000000000010001101001111",
"00101001011010000001001110011010",
"01010101100011010011000111011101",
"10110110100111010111011001000011",
"11001000010100000001100111011111",
"10001001001101000010000100111110",
"11110101101101011110100111001000",
"01100000000011010101111100110010",
"00011110111001111100100100101111",
"01011001110110111001100100111110",
"00100101000101010011011110111100",
"01001100101110111001100001010011",
"00110010001011101010110010010101",
"01111001000101101000000101110111",
"00000101110110011011100000100100",
"00111110110110001000010001100001",
"01000000000101110101011101100101",
"01110111101110010111101010001011",
"00000111001100001010101011001110",
"01001110101110101011111000101000",
"00110000001011110111100010100111",
"00100011100001111101010111010011",
"01011011011100010011101111000000",
"11011001111000100110000010100011",
"10100101000100001011111111010111",
"00010011001110110000101111101000",
"01101011101011110010111110110110",
"01110011000100001111011000010010",
"00001011111000100000101111110011",
"01001110010010101000010101001101",
"00110000101000011100110011111101",
"01001101100111011001010100010010",
"00110001010011111111000100101111",
"10010111100010101000101010000011",
"11100111011011001000010110011110",
"01110010010011110011100001001001",
"00001100100111100010000110101110",
"10110011000000101111110000111111",
"11001011111110100010101001011000",
"11001001000011111010010000001100",
"10110101111001000001111111100101",
"10000101000000011110110101100000",
"11111001111111000011001111100011",
"11001110000001100100011010110110",
"10110000111101000000100011000111",
"11011110100100011101100110011011",
"10100000011000001010101101001101",
"10000010100101000011001011111011",
"11111100010111010001101110011111",
"10110110111111010101101010001011",
"11001000000000010101011001000100",
"01101011000101010000110110000111",
"00010011110110111101011101101100",
"10011000001000011111101010011001",
"11100110110010100100110001000111",
"00011100100110110011110001110111",
"01100010010100110001010110110101",
"10111010001111011111011101100001",
"11000100101011000111111001100101",
"10000100100101111100101111100000",
"11111010010101111101111000111101",
"00101100001001010011110000110101",
"01010010110001100100111110110000",
"10001101011100000111100000111111",
"11110001100010000100010001000011",
"10011111001101101010001001110110",
"11011111101100110110101100011001",
"11100100011011100111001001111011",
"10011010100010010110110000100111",
"11010010000111000100100000000100",
"10101100110100011010110001010110",
"01011111000110000011010000110010",
"00011111110101110100101001001000",
"01000011010010010101001011100111",
"00111011101000101100001100111101",
"01010101001101101010010000111011",
"00101001101100110110100101011100",
"00111001111111010100011000000000",
"01000101000000010110000011000010",
"11111000001001101000000010101001",
"10000110110001001100110101000000",
"10101001000110011100100001011001",
"11010101110101010001010001111100",
"11001011011111111101000011101010",
"10110011100000000001011110001111",
"10101000001100101111110001011100",
"11010110101101110001001101110101",
"11101100100110001100100101110101",
"10010010010101100111011111110110",
"11110111110001110011111111101011",
"10000111001001000111010011111100",
"01101010111110010111000001101100",
"00010100000000110101110111100001",
"01000011011001011111011001000111",
"00111011100011100111111000111011",
"11100111100111000100001011011001",
"10010111010100011011001101000101",
"01111000001010011001100100110101",
"00000110110000010011010110010100",
"10110100110101100011011101110010",
"11001010000110001111011101111000",
"11111001100010001100101111011100",
"10000101011011111000100111100010",
"10100001011001000001011010011110",
"11011101100011111010100111100100",
"11000001000011001110011010001101",
"10111101111010001000111110100110",
"11011110101011010100101101000101",
"10100000001111010001011011001011",
"11001110011001011001001000010000",
"10110000100011101011110001101111",
"11101100000001001100110100011001",
"10010010111101101011111010101101",
"10111010000011110101101000100000",
"11000100111001001001010110001000",
"00111000101110110001110101011100",
"01000110001011110001111101011111",
"10011111100111111010101101100100",
"11011111010011010011100101010011",
"11000100101100110100101000111001",
"10111010001101101100001111110011",
"00010110100001000111110000100110",
"01101000011101110101010101110000",
"00111011010100110110011101110000",
"01000011100110110000000001110011",
"10101000000101101010001101010010",
"11010110110110011000011100110101",
"10111100100001110000101100101011",
"11000010011100101010010111000100",
"01101110111110100101111110011110",
"00010000000000101110000001100000",
"01101010100001100001110111000000",
"00010100011101000101001101001111",
"00000101010010111010111001000011",
"01111001101000001110000100010111",
"00100101010101010100101000111101",
"01011001100110011010000110010111",
"00000010100001001110111100111000",
"01111100011101100111111101011000",
"01000001011000101100000101011110",
"00111101100100001000001000011000",
"11011010110101100110000101110001",
"10100100000110001101100110000001",
"11001000011010011101101110110001",
"10110110100011000001111001111110",
"01100100111011000010110001111010",
"00011010000010101011111011001101",
"01110111001010000001001000001101",
"00000111110000101111011100111110",
"10100110011110001101111111011111",
"11011000100000111010101000101101",
"00011011111100101100001100101110",
"01100011000001101111101011001110",
"01101011100010000001011011101101",
"00010011011100001100100001011010",
"10010110111001111100111001110100",
"11101000000011010101101111111011",
"11111010001101011101010011100111",
"10000100101101000011010111101101",
"10110011110111101111011011000110",
"11001011000100101111011100101000",
"01000100110011000001110000111101",
"00111010001000001000101001101000",
"01010001101100110101111111111111",
"00101101001101101010110111000011",
"00101010010011110100100011100101",
"01010100100111100001010100000010",
"10010000011100000101111101010001",
"11101110100010000101001001100101",
"11111011000010110011111110111111",
"10000011111010110101000111000111",
"01111101101111101011100101100101",
"00000001001010111100111011101101",
"01101010110001110101110011000010",
"00010100001001000101110100110010",
"11000111010011011000111000100100",
"10110111100111110110100110000010",
"01101000101100101011001101111110",
"00010110001101110101111000011011",
"00011101110010101100101100010110",
"01100001001000011001010101001111",
"10101010110000111100101000001010",
"11010100001001110101110100011001",
"01011011111010111010000101001010",
"00100011000010110001000011000010",
"00011100111100011001110001000010",
"01100010000001111001111110010001",
"00010101000110100111001000011101",
"01101001110101000010101001000100",
"10111111010100011010101010110111",
"10111111100111000100100100111001",
"11101111001101011010011110001111",
"10001111101101000110001011101001",
"00100011111111100101100011011011",
"01011011000000001101010011110010",
"00001000000011011011010011110011",
"01110110111001110011110011101011",
"01000110010110010010100010010001",
"00111000100101101110010011111001",
"00000110010000011101100011011011",
"01111000101010010000101001011011",
"11011000111110101001010111100011",
"10100110000000101100010000001000",
"10001010010000000111011100001100",
"11110100101010100100000100011010",
"11101001101000110110001110100001",
"10010101010010001000110101000101",
"00100101101100010110000101110100",
"01011001001110001011101110001110",
"10111111010101000111001100110101",
"10111111100110100011110100010110",
"11010110111110111000110111001100",
"10101000000000100100001100101001",
"11001100110011110000111010001110",
"10110010000111100100000110001101",
"10101011110000111101010110111101",
"11010011001001110101001100011001",
"00001001000010001010010101001001",
"01110101111011111100110110000000",
"00111010100100010011110111011001",
"01000100011000011001110000111101",
"00011010110001001101011000110101",
"01100100001001100111100100010101",
"11011001010111110101101010110111",
"10100101100100101011010101100101",
"11000011010010111101010111011100",
"10111011101000001100000111010110",
"11110011001100011110011100111101",
"10001011101110000011000010100010",
"11100100100001100000010001011101",
"10011010011101001000000110010111",
"01001101101111001110000001100011",
"00110001001011010111110100110000",
"00000001010000101000110011100101",
"01111101101010000110110111101100",
"00101001100010110101110010100001",
"01010101011010110010000100000010",
"00111010111010011100001011011100",
"01000100000011000010110101100001",
"01101010011100000001101011100101",
"00010100100010000111100100111101",
"11010010111110000000110100010101",
"10101100000001000001101000010000",
"01000100110011000111111110111111",
"00111010001000000011110001001001",
"00100000111111111101010001000100",
"01011110000000000001010111100010",
"00111111100110100010101010101100",
"00111111010101001000110010010110",
"00010110001011110111010100001001",
"01101000101110101100001000000001",
"00000101010101111111011110000110",
"01111001100101111011101000011010",
"10011001001000100010111111110011",
"11100101110010100000100110111011",
"01010000111110111101111101101011",
"00101110000000100001100011110011",
"11010010010010001100101111010000",
"10101100101000110011000010111101",
"00000101110001111101011101001001",
"01111001001000111111100001101100",
"01110011000000100111111000001001",
"00001011111110110001110001001101",
"11111000000000110000001110100100",
"10000110111110100001110000111010",
"11101101010010111100101100100000",
"10010001101000001100101001001110",
"00011011001110001111100101001001",
"01100011101100010010011001000010",
"00001010011011100011000000011011",
"01110100100010011001001001110010",
"00111010000110101101111010100100",
"01000100110100111001010110010111",
"00111100111010000011110110100001",
"01000010000011010001100001010000",
"01011100001000100010000000000010",
"00100010110010100001110110011001",
"01001100101111001000001101101100",
"00110010001011011101001010111110",
"10111001011110010010010000000100",
"11000101100000111000011000101010",
"01110110000110110100101110010000",
"00001000110100110000000100110000",
"11010010011110101100100000110110",
"10101100100000101010100111001011",
"10000111011101001110100011101101",
"11110111100001011100101111010001",
"00011011100100011001001010110100",
"01100011011000010001100010111010",
"11011000111110001000101101101010",
"10100110000000111101011011101011",
"01111001110000110110000011110010",
"00000101001001111011011100011111",
"00100110000100011000100101100001",
"01011000111000010010011100100110",
"11000000010000000001010001100011",
"10111110101010101001100010001101",
"00010011010101001100010011011011",
"01101011100110100000000111100110",
"00111011100100101110001001111101",
"01000011010111110001011000100110",
"01100001001000100010000111011010",
"00011101110010100001101101001100",
"11111011001010010011001000100110",
"10000011110000011010101101000100",
"01110100100101010001111110000110",
"00001010010110111011110011100101",
"01111011111100100111000101100001",
"00000011000001110010100001011001",
"11110011000001111001110011010110",
"10001011111100011010000100100000",
"10100100001111011001101101101000",
"11011010101011001101001000010001",
"01110100001111001011000011110000",
"00001010101011011010100011010001",
"11111000011000000110001111101010",
"10000110100100100000100000000010",
"00011010001011110000101100111111",
"01100100101110110011001011011111",
"01010101011011110100111010011011",
"00101001100010001110110110111110",
"10110101010010110110000010011100",
"11001001101000010001111010000100",
"10111111001000101010000000011110",
"10111111110010010111111001100001",
"11000000111110010001010000100011",
"10111110000000111000111010001101",
"01101110101110100011111001111111",
"00010000001011111111000011101101",
"01011010110110111100001000101101",
"00100100000101010001101111110000",
"11110010000100001100110111110100",
"10001100111000100100101010010011",
"00011111111110101110001000011110",
"01011111000000101001110001001101",
"01011010000010000100001110000010",
"00100100111100000111100110010011",
"01000100100001010101001001000010",
"00111010011101011100100000111011",
"11010101111000011010010010010111",
"10101001000100010011100001111001",
"10001011011001100100101001001001",
"11110011100011100100101001000001",
"10100000101011111101011110000000",
"11011110001110100101100101101101",
"01110000110101111010001110011101",
"00001110000101111111010100100101",
"01111011010101001001010100010111",
"00000011100110100010010010000001",
"00101101000000100011001000001001",
"01010001111110111010111011100010",
"11111110001011100100010110000110",
"10000000101111000000011101000011",
"00011111111101101001001101000000",
"01011111000001001110010001111100",
"10111101101010100111110010100010",
"11000001010000000011001111011000",
"10111100101100111001101000100101",
"11000010001101100111001010011110",
"00110101001111011000000001100010",
"01001001101011001110101010110110",
"01010110101100011101110000011110",
"00101000001110000011110000100111",
"01010011100011010100000001011001",
"00101011011001111111101111001110",
"00010100100010000100111001110001",
"01101010011100000110011001001001",
"10001011001111001011111111100001",
"11110011101011011001101100010001",
"00000011100100000011100011000000",
"01111011011000110011010010101110",
"10010000100110101000111111001100",
"11101110010101000000000110000101",
"01011011001111011010010001110111",
"00100011101011001100100111010000",
"00001110100110010111111001000011",
"01110000010101010111101101010100",
"01001010010110101010001010110111",
"00110100100101011101111111111101",
"01010111000110111111011011110000",
"00100111110100100001100101010101",
"11011010101100011111011100001100",
"10100100001110000010000001000110",
"01011001101010100110011101100101",
"00100101010000000100101111001100",
"10010010100110110010001000011011",
"11101100010100110011100110010011",
"11011011100110000011000110110000",
"10100011010101110100110111010100",
"01000011101110011001111100101001",
"00111011001100001000011111110100",
"11100110110111100001100010010011",
"10011000000100111000101000110001",
"10111000001001000000000001101000",
"11000110110001111100110110001110",
"10010001000110000011100110000011",
"11101101110101110100001011000011",
"01101000000000001101110011001001",
"00010110111111100100100101100011",
"10100101101110011110111110001101",
"11011001001100000011101110100001",
"11111101011100110101110111011100",
"10000001100001101010010100000100",
"11111010100001111001100010010010",
"10000100011100011010100010111010",
"11100111100111101110011010100110",
"10010111010011100011011101101100",
"10100100110001100100101001100111",
"11011010001001010100000010011100",
"00010011000011110010101000101111",
"01101011111001001110001000010011",
"00101001010101100101111000011101",
"01010101100110001101101111100001",
"01010001001011000111110111001111",
"00101101101111011111100000000110",
"01101000011010011010101110001000",
"00010110100011000011101101011111",
"00011010010101011010100110001001",
"01100100100110010101110100010001",
"00110011000101100101110000101011",
"01001011110110011110111000100101",
"11010100110101111000111101001010",
"10101010000110000000001101111000",
"11111000011110101100001111111001",
"10000110100000101010110000000000",
"11010100010111111100110110101100",
"10101010100100100110101000001010",
"11011001101001111101111010001100",
"10100101010000110011001100001111",
"10100101111001111111011011100001",
"11011001000011010100001101011001",
"00100111111100011011111111111110",
"01010111000001111000101110000101",
"00110101101101100100110101110011",
"01001001001100111011111011000011",
"11111100000011000101011100010001",
"10000010111010010111110101101100",
"10101011100110100110111101100110",
"11010011010101000010110111111111",
"11001111010011101011110101110110",
"10101111100111100111111110100000",
"10011100101101001110001011010001",
"11100010001101010010011100011100",
"00101100011010101011101011010001",
"01010010100010111001100101001101",
"01111011101001011110000100010101",
"00000011010001011000101010010011",
"01010001101010010000000010001010",
"00101101010000011110010000011110",
"01011000110101100100001110010010",
"00100110000110001110111011010000",
"11110100000010101101001101010001",
"10001010111011000000100110010011",
"00011110101100111101000101110101",
"01100000001101100011101001111111",
"10111010101010010110001010010000",
"11000100010000010111001111101001",
"01110110000110001001010011000111",
"00001000110101101100001000000010",
"10101111011101000100100110010110",
"11001111100001100010001100010110",
"00010011101100110000111100110110",
"01101011001101110000000000101110",
"10111111010110111110000001100111",
"10111111100101010000011101110001",
"01111001110111110110001000100100",
"00000101000100101011000010000101",
"01100110101111101001000011000010",
"00011000001010111111001110010000",
"01011100001110101101100011110001",
"00100010101011110101111101111111",
"01100100001000110110101100100000",
"00011010110010001000010000010010",
"10101110101100100110100111001011",
"11010000001101111010100111011010",
"01100110110100010001110001100010",
"00011000000111001011001110011010",
"10100101011000101000110001001011",
"11011001100100001010001111110010",
"01000000010100111101010101111110",
"00111110100110101010111111101100",
"10111101001110010111100110100011",
"11000001101100001010101110101011",
"00101011111001101010001010111011",
"01010011000011100001001110110000",
"10100000111001000100000000011010",
"11011110000011111000111111000111",
"11001111000000001110101000111001",
"10101111111111100010111011100001",
"11111010111000010100011001100111",
"10000100000100010111010100110000",
"10110010111111010110000010001010",
"11001100000000010101001100110101",
"11010101110110110011110101100011",
"10101001000101010111011001000000",
"11010111111111011011001001000110",
"10100111000000010010100110001010",
"00101101110000010111100001101010",
"01010001001010010101111010011111",
"11110101001101000111000100010010",
"10001001101101011001100101001110",
"01110100110010011001000101000000",
"00001010001000101001000011100100",
"10000010111011000000110100011110",
"11111100000010101101000100111100",
"01101001111001100000001000100011",
"00010101000011100111011011100011",
"11001101110101000100010111101011",
"10110001000110100101110111111111",
"00100010001101110100011001101101",
"01011100101100101100101010010101",
"00001101100000010101111001001101",
"01110001011111010100101011001111",
"01000010100001101100010000111001",
"00111100011100110010010110000000",
"10111011010111100000101100101000",
"11000011100100111001001100011011",
"10011111111110000000011001010011",
"11011111000001000001110110101010",
"01111010011001111101100100110101",
"00000100100011010101010101101101",
"10001000110101000010100100110000",
"11110110000110100111001011100110",
"10101001011011011010001001011000",
"11010101100010011110010010000100",
"00011111101111100111101010110001",
"01011111001011000000011101111011",
"10101110011010100000011000011011",
"11010000100011000000010100011001",
"11000000001001111001011110100111",
"10111110110000111000010110100010",
"11010111011111000100010001110110",
"10100111100000011110010011010111",
"01111100111101100101001101011111",
"00000010000001010000011011110011",
"01011000011011010010001111110011",
"00100110100010100010111000000011",
"01000100001001010111101100010101",
"00111010110001100000010001010110",
"01110110001001001110001111110001",
"00001000110001101011100111011000",
"00110100011010011000010101001000",
"01001010100011000101001001011000",
"01000101110011011000000110010011",
"00111001000111110111001101000001",
"10111101000011100100001101000110",
"11000001111001100101010110010101",
"11011010010110110100110111010101",
"10100100100101010110101100001011",
"00001011100010101000001000011101",
"01110011011011001001001111110101",
"11110111110111111001011001010100",
"10000111000100101000111001001000",
"00000010001010000110000011001010",
"01111100110000101001110000010010",
"11110011000011100001000111100001",
"10001011111001101010010110101010",
"00100010101110001000110101001010",
"01011100001100011000110111101100",
"11101111011001101100111010010110",
"10001111100011011111100010110001",
"01000101000101101000111100101001",
"00111001110110011010010001010110",
"00010111110100010100110111011001",
"01100111000111001000111010010001",
"00100001010010110110010010100001",
"01011101101000010001101101010100",
"00101000111010010011100000001010",
"01010110000011001000000011010001",
"00010110011111111101101110101010",
"01101000100000000001001000101110",
"11001011110011011010000100111000",
"10110011000111110101101010111000",
"10100010101101000101111000111010",
"11011100001101011010110001000111",
"11000001110110011010101001110101",
"10111101000101101000101011101101",
"00010010110001101010111110000111",
"01101100001001001110110010000000",
"00111100110010001110101100011010",
"01000010001000110001011101010011",
"01110000111110000001111101010101",
"00001110000001000001000001011001",
"10110010101011111101110011110001",
"11001100001110100101001110101001",
"01010101111101011011101000011010",
"00101001000001010101100111101100",
"10010101000001110101101110011010",
"11101001111100100001010110010011",
"01000111001101100000011011001110",
"00110111101101000000010010000110",
"11011011100011100110110001010110",
"10100011011001100001001100101100",
"11001011010100010011110100111100",
"10110011100111001001101011111111",
"11001110010110010111100001111111",
"10110000100101101010110110000011",
"01100011100111100010101111111011",
"00011011010011110010101011001010",
"01010010000011011000000110010011",
"00101100111001111001000011011111",
"00010110010100001100110010000110",
"01101000100111001110111110001001",
"01000101000001110110100010011001",
"00111001111100011111111001010111",
"00101111011101100100010110010111",
"01001111100001010000111001100101",
"00011000110001111100110001000001",
"01100110001001000000000101111001",
"00100011000101100000101101011000",
"01011011110110100110001110001010",
"11100000100011100010011011000010",
"10011110011001101000001111001001",
"00001010001110010011100011001010",
"01110100101100001110100110000101",
"10000111001011101010101011001100",
"11110111101110111001101000111110",
"00111000111110111111001010000110",
"01000110000000100000111100010101",
"11011000110111010011101001001010",
"10100110000101000001111001110000",
"00100000101001000011000010010110",
"01011110010001111001001011101101",
"10001100011111101000111101001100",
"11110010100000001011100101100101",
"00100111110010110110000011010000",
"01010111001000010001111001011010",
"11011000100100100000111110110000",
"10100110011000000101100000011101",
"01010010000110101011100001010110",
"00101100110100111100100111111001",
"00000101100001111001010001110001",
"01111001011100011011000000010110",
"01001000011110101011010000010000",
"00110110100000101011010001001011",
"10100001011100001010111110011100",
"11011101100010000010010011101010",
"01010001011100000001000000011000",
"00101101100010000111111101100001",
"10111010001011011110111011000110",
"11000100101111000110010100001011",
"00001111110010010011001100111010",
"01101111001000101101110011011100",
"00001000100101000100011000011110",
"01110110010111001111111100010101",
"10101101111110100001100100111100",
"11010001000000110000010100110101",
"11111010001100010101111011101001",
"10000100101110001011111000110100",
"10101011111110001111011101010001",
"11010011000000111001110111000111",
"01100111001010000000010100011000",
"00010111110000110000011001000111",
"00000111011110100011111111010100",
"01110111100000101111000100000000",
"00111000100100101001010110111011",
"01000110010111111000101011110111",
"11001110011111101001110000110000",
"10110000100000001011001011100001",
"00111010101011110010110101101111",
"01000100001110110000111001010111",
"10111011110001000011011010101111",
"11000011001001110000000001101101",
"10001001000001001101100101100010",
"11110101111101101010011111011100",
"10001010110001011011111011101011",
"11110100001001011011010100101101",
"01111100001011111110010001100111",
"00000010101110100100101111000010",
"11100100101011100000010011011101",
"10011010001111000100110100100001",
"11010000101110111110101001110101",
"10101110001011100110000000111101",
"11010001000110011110100010110101",
"10101101110101001110011110101111",
"00001110011110011010010000011011",
"01110000100000110100001010101110",
"11101001000100110010000101111110",
"10010101110111101011011010011110",
"01100110000010100000110110110101",
"00011000111011010101101101110000",
"11011011101110011001110000111000",
"10100011001100001000101011000000",
"01100001101010010100000010111000",
"00011101010000011001101010011000",
"11000000110110001010011100110001",
"10111110000101110011111100010100",
"00010010011110010111110010110000",
"01101100100000110101011101101011",
"00101011011000000111101111011110",
"01010011100100011111100001101101",
"00101111111100001001011111101000",
"01001111000010000011001001010100",
"10001101010111110110110000000001",
"11110001100100101010101000001011",
"01101011011000111001110101001101",
"00010011100011111111011001110110",
"01100011011010101111101001001010",
"00011011100010110111001110011000",
"11110100010110101111100111110000",
"10001010100101011010010001001010",
"10011101111100010101010011100001",
"11100001000001111100011110101110",
"10111100100100000011011100111110",
"11000010011000110011011100001110",
"10011110011001110001010011111001",
"11100000100011011100110101110010",
"11101110000111110011111110001001",
"10010000110011011100010001010001",
"01010011101101001101111001011110",
"00101011001101010010101110010001",
"10011100100001100100111101000111",
"11100010011100111111100100110110",
"10100001010110110110000000001011",
"11011101100101010101111010100100",
"00010010101000100101011010100011",
"01101100010010011101100110010101",
"00011000011010110110011001110010",
"01100110100010110011001110000101",
"11110001100010110100101010011110",
"10001101011010110011111101101010",
"11110010010001000111110101110100",
"10001100101001101100010001000111",
"10101010111100001001010011011111",
"11010100000010000011010000001100",
"01011010011100010101001111010010",
"00100100100001111100100001000111",
"00010111110010010001010001100001",
"01100111001000101111010111011001",
"01111101111001111011001111100001",
"00000001000011010110110000110010",
"00000101111101010100110101000011",
"01111001000001011001010100010111",
"11010001001110101111001010110111",
"10101101101011110100011101010010",
"00001010111001000100011001011001",
"01110100000011111000101111011010",
"00001101100011110101111111011010",
"01110001011001001000110001100111",
"11110111000111000011111000101000",
"10000111110100011011100110010001",
"11001101001011001101001100100000",
"10110001101111011001101000111111",
"10010000101100101011100011010000",
"11101110001101110101100010100110",
"10010001110100100001110101101111",
"11101101000110111111001111100101",
"11010000101111000011101001101000",
"10101110001011100001011000101100",
"01001000011100001110001011000111",
"00110110100010000000011111111111",
"11101110000010010110011000110010",
"10010000111011100111110011010001",
"11100011110000110110011110001101",
"10011011001001111011000101110100",
"10111010010110010100100110110000",
"11000100100101101100110111111000",
"00101111010011100010110100111110",
"01001111100111101110111001111110",
"11111100000100010000100101111011",
"10000010111000011110110110110010",
"01011110010001100110110001100100",
"00100000101001010010010001001110",
"11001001000011101110100111100001",
"10110101111001010100100100010000",
"11000100100010111101101100111111",
"10111010011010100100110000100011",
"00011111001000110110011011001100",
"01011111110010001000100101100010",
"01001100111101101011011000011101",
"00110010000001001101000110110101",
"00110011010111110111100101010011",
"01001011100100101010000101001101",
"10101001111000100011001001100011",
"11010101000100001101110101110000",
"00001000101010111011110001101001",
"01110110001111101100110111110101",
"11100111011001110100000110010110",
"10010111100011011011001000010111",
"01100101111100011101001110110100",
"00011001000001111000000001111001",
"00011011101011110111101111011000",
"01100011001110101011101011000010",
"11101010100011011000010010011001",
"10010100011001111000101111101101",
"01101100111101010011010011111000",
"00010010000001011010001001010011",
"00111101101001111001111011000101",
"01000001010000110111110101010101",
"01110111000010010010110001011100",
"00000111111011101110000101011110",
"01001001011110010100001101010101",
"00110101100000110111010110100100",
"00111011101111101111111011111111",
"01000011001010111001000001010001",
"00000100110100001111011111011011",
"01111010000111001100111011111110",
"11100110011110110101110101110001",
"10011000100000100101110000111000",
"11010010011001100001010101011000",
"10101100100011100110101011111110",
"10111010001101000000001110011011",
"11000100101101100000011110111011",
"11001101100101011001110011001101",
"10110001010110110000010011100110",
"01001001110101111100000011001110",
"00110101000101111110000010010101",
"10011111110010101000010111010001",
"11011111001000011100110010010100",
"10101111101010010101000000001000",
"11001111010000011000100100010101",
"01100001000101110010011011000011",
"00011101110110001100101000001100",
"01011001101101111001001101101100",
"00100101001100100111111110011000",
"01001010110010111010111101000101",
"00110100001000001110000001001011",
"01110000100010110111100110100110",
"00001110011010101111000000010110",
"01100010111100000010101010011010",
"00011100000010000111000001010001",
"11000010001010111111011001001011",
"10111100101111101000110110111011",
"00111100111001000011111011000010",
"01000010000011111001000010100000",
"00111110111100011001101100100101",
"01000000000001111010000000110001",
"11111110001101011100111110001000",
"10000000101101000011101101000000",
"11100101101010011001010101000101",
"10011001010000010011101000010001",
"11011000110111110000110000100110",
"10100110000100101110100100010011",
"11010110011000010111001110001100",
"10101000100100010101100000010000",
"10000011111100111100111011100000",
"11111011000001100110011010011010",
"11111100101101100000001000101001",
"10000010001101000000100100011110",
"11010001011110000011011011000000",
"10101101100001000000001111100011",
"10101001011110101010111000110111",
"11010101100000101011011101010111",
"11110111101110000001111000010001",
"10000111001100011111100100101110",
"11111110001101000000100011011111",
"10000000101101100000001001101000",
"01001001110111110000101000000111",
"00110101000100101110101001111000",
"11001010111101110001101101100001",
"10110100000001001001101101000111",
"01010110010101000010100010001000",
"00101000100110100111001101100001",
"11011001001110001010001010010000",
"10100101101100010111100101110111",
"10001011000011100000011011110110",
"11110011111001101011011101100101",
"11010100111011011001110111101001",
"10101010000010011110011100010110",
"00111101100101110011011001001100",
"01000001010110001011001111000110",
"01011001110111111011101101100000",
"00100101000100100111011000000011",
"01011010011101001100110000001111",
"00100100100001011101101110011000",
"10111100111010101110101101100101",
"11000010000010110111110001101111",
"11010000011110100110001101000111",
"10101110100000101101111001110110",
"10000010001001101110111110100001",
"11111100110001000100101001101110",
"01100110000000000011111111000000",
"00011000111111111000000010111111",
"01010100100000011111011110001010",
"00101010011111000010000000101010",
"00101110110100111101111101111011",
"01010000000110101010100010100001",
"00100000001111000010101100101001",
"01011110101011100010010001000111",
"01000001011101011000001011110000",
"00111101100001010111011111100011",
"00100101100000100001111000100011",
"01011001011110111101010101100000",
"11111000010101100101100000110111",
"10000110100110001110000000010110",
"10101011000000100001001011000011",
"11010011111110111110101101100110",
"00010110111001001111111001101000",
"01101000000011110001100001111001",
"10001100101010000011010110101100",
"11110010010000101100110111110101",
"00111010100001101110001111011011",
"01000100011100101110110001111011",
"01101010111100100111011100100111",
"00010100000001110010010100100001",
"10010110110010010001111111111001",
"11101000001000101110110001110100",
"01110011011001000100101011011010",
"00001011100011111000100100000101",
"11100001011111100101000000011100",
"10011101100000001101100101100001",
"00001001001101100001110101001000",
"01110101101100111110111001001110",
"00100001001011001101100001010011",
"01011101101111011001010010001011",
"00100101001101101110110110101110",
"01011001101100110010000101010010",
"10110000011011100001010100111100",
"11001110100010011010000111111001",
"01001000101100111010000101010000",
"00110110001101100110101101010111",
"10110000101001100101111101100010",
"11001110010001001111010010011101",
"10001001101011010100001110100101",
"11110101001111010001111100011110",
"01101100111100001000000000100110",
"00010010000010000011111111001000",
"00101100011000010001011011000110",
"01010010100100011001001111111000",
"10110100100111110000011100010101",
"11001010010011100000110101011101",
"01011000010100011011001101000011",
"00100110100111000100001011011010",
"10011111100100010011110101111111",
"11011111011000011001110011001001",
"00000100001000011001101011011010",
"01111010110010101100010000100010",
"01101011001000011000110011111000",
"00010011110010101101010110001111",
"00011101100111011110000010111001",
"01100001010011111000110110001011",
"11101101000100010010000000101111",
"10010001111000011100101001011010",
"00010100000111100110110011110000",
"01101010110011101101010111011001",
"10000100100011000001001011010011",
"11111010011010011110111100101101",
"01011110001111101011000001010000",
"00100000101010111101011100011100",
"00100110110111011100000000111100",
"01011000000100111100010011110111",
"10010101001010000001000100010011",
"11101001110000101111100001100000",
"11011000011010111000101001110001",
"10100110100010110001111000111111",
"01100101001110100101101001001010",
"00011001101011111101011010110000",
"10000101111011100000111111001000",
"11111001000010011010010100100000",
"10111101110101011110110110101011",
"11000001000110010010110000111001",
"00001000111111110100110001001111",
"01110110000000000101101000011000",
"10100001100000111110110101110110",
"11011101011110000110000011110010",
"00010011110000011000100010100011",
"01101011001010010101000001101100",
"00000100101001101100110011011110",
"01111010010001000111001101010110",
"11011001010001010101011110000010",
"10100101101001100000110000000010",
"11011000001100110110011101011101",
"10100110101101101010011001000011",
"00100110101110010001111100010010",
"01011000001100010000001000011001",
"00010001101110011010001001000000",
"01101101001100001000010100000100",
"10000101001001101110011110000001",
"11111001110001000101001111111100",
"01010100111100000110010101100001",
"00101010000010000100111011110100",
"01101001001000100110011001011110",
"00010101110010011100011000001000",
"00011100011001111000100111001110",
"01100010100011011000010111100101",
"00110010001010001001000100001010",
"01001100110000100110010001011110",
"11101000001101100010001000000111",
"10010110101100111110100110011110",
"00000000100101010101110010100001",
"01111110010110110110001011111111",
"01001101011001011010100111100000",
"00110001100011101010110110100011",
"11111110010101100101010110000000",
"10000000100110001110001000000101",
"00101110101111101100010010000110",
"01010000001010111100010011100111",
"10010010100001101001101111011111",
"11101100011100110110111001100100",
"01110100101101010000111101101011",
"00001010001101001111101001111100",
"11110101011001111110000001111100",
"10001001100011010101000011111101",
"01000111011110010111110101101100",
"00110111100000110101011100001000",
"11010010110111111000101011011100",
"10101100000100101001010111001101",
"11000001101000101001001000010110",
"10111101010010011000111111000101",
"10010001110010101000001000101010",
"11101101001000011100111101111111",
"01110010010101010110101011110001",
"00001100100110011000101000001100",
"11000011111011101110011101001010",
"10111011000010010010100011110110",
"01001001010010011010100100110001",
"00110101101000100111110110011000",
"00110001000100101000111001010101",
"01001101110111111001011001000000",
"11100110000101011111011100001010",
"10011000110110101000000100011011",
"00100010101101010011100110001111",
"01011100001101001101000001100111",
"11010011110000010011010100001111",
"10101011001010011001100110101010",
"10010100101000101101001101101101",
"11101010010010010011111011100011",
"00100100000010001011000101101101",
"01011010111011111011100000110100",
"00001010100001000001010110011110",
"01110100011110000001010101101111",
"00010001111000110111001010001000",
"01101101000100000001000110001000",
"00001101011010001011010111010100",
"01110001100011001100111101101111",
"00011100000011001111010110101000",
"01100010111010000111011010111010",
"10110010100100000000111110100001",
"11001100011000110111010110001001",
"10111000010011101011001100001101",
"11000110100111101000011110011100",
"01110100010000100111111100110110",
"00001010101010000111100111000110",
"00111111010001110111101001010100",
"00111111101001000100010011010101",
"10111001011000010001001010111110",
"11000101100100011001011010010011",
"10101110010010001101111011010101",
"11010000101000110010000101001001",
"10111010000100001110111010111101",
"11000100111000100001011101100010",
"00011100000110111000110000001010",
"01100010110100101010100110111001",
"11000111110110100111011011001001",
"10110111000101011111111000100000",
"01111101110100011011011101011011",
"00000001000111000011111111001110",
"01110010010111001011101010101111",
"00001100100101000111010000010001",
"10000011101001101011100110000010",
"11111011010001001000101000100110",
"00111010100110000010100110100001",
"01000100010101110101100100111011",
"11111100110011001100011001101000",
"10000010001000000000010011111111",
"01101110111001110001101111111110",
"00010000000011011100100100100100",
"00101000010010010010000000100101",
"01010110101000101110110001010000",
"01110110100010010100001111001111",
"00001000011011101011100010001111",
"01100101110100011011110101101011",
"00011001000111000011101101001001",
"10001011001110111111000100110000",
"11110011101011100101100111111110",
"00100010111111010010100110000110",
"01011100000000010110111101001111",
"10101101101010100101101101000100",
"11010001010000000101100101111101",
"00101111000100001010010100000010",
"01001111111000101000101010100010",
"01100101101001001101111000111010",
"00011001010001101100000010111011",
"11000100100000010111001001001110",
"10111010011111010010001110101011",
"00111011000010001111001000100110",
"01000011111011110100011011101000",
"10001001111111001001111100111001",
"11110101000000011011011000101100",
"11100100001011011001001001110010",
"10011010101111001100100101000001",
"10101010010001100111110100100010",
"11010100101001010001011001100000",
"00100011001011011000010011000101",
"01011011101111001101100000100010",
"01100110110001101001101110001000",
"00011000001001001111110100011011",
"10111111111011001111111110011011",
"10111111000010100100001100110011",
"00110011100010111100110001100100",
"01001011011010100110010100001001",
"11101111101001111000111011011111",
"10001111010000111000111111100001",
"00100001010000100000011001110000",
"01011101101010001110001010100101",
"10111110011101101100000110001111",
"11000000100001001100101110001100",
"10111111100000001000001111111110",
"10111111011111101111100100010011",
"00010101100001010011100001010010",
"01101001011101011111100000010101",
"11010011110111000110011011010101",
"10101011000101001010110010001011",
"00111001101111010101101000001101",
"01000101001011010000110110110111",
"10101000101010010110101110010000",
"11010110010000010110100110100010",
"01011010101100010000001011001110",
"00100100001110010001111001010101",
"00100010001010111111100100001000",
"01011100101111101000101010110010",
"01000000010010010110001110000101",
"00111110101000101011010111001111",
"11011101101001000101000101010100",
"10100001010001110110101100101000",
"01110011100001011011100110110101",
"00001011011101010000101000011000",
"01110101100010111000100100001111",
"00001001011010101101011000100100",
"11010011011110101010100010001010",
"10101011100000101011101001001101",
"11101001111010001111110010111010",
"10010101000011001010010010010110",
"11000010011101001101111101000010",
"10111100100001011101000100011010",
"10111110000001011011011101111001",
"11000000111101010000111000110000",
"01001111011010100011001100100010",
"00101111100010111110101000101110",
"01101101000011001011110110100101",
"00010001111010001101001100111110",
"01101100000101110110010001111000",
"00010010110110000111000110101111",
"11100000000110011000001000000001",
"10011110110101010111011000100000",
"01011001010001101111110110011110",
"00100101101001001010101111001000",
"00011010100110110000101010111000",
"01100100010100110101100101110000",
"00111011011010001111100001011100",
"01000011100011001010011100111001",
"11110010110101101001010110101101",
"10001100000110001011010001001100",
"10001001001110010111100111101011",
"11110101101100001010101101100110",
"01011111001010010100010000101100",
"00011111110000011001011010100101",
"10010100111001011101001111011101",
"11101010000011101001001110010010",
"10110000001100011110110011110000",
"11001110101110000010101010111100",
"01111101110011000010001010101110",
"00000001001000001000010101010111",
"10101011100000101011001111010001",
"11010011011110101011010011111010",
"00100101010001011110110011010101",
"01011001101001011000111010111100",
"11000001001011001010001011000010",
"10111101101111011100111101011110",
"11100111000011101010011011000010",
"10010111111001011011010011110011",
"11011001100111111000101101101100",
"10100101010011010110001001110010",
"11101111001000101000010011100010",
"10001111110010011010000000100101",
"01111000111110101100100111000000",
"00000110000000101010100011111101",
"11000010011110111111101011111111",
"10111100100000100000101010110110",
"11111100011000011000001011101101",
"10000010100100010100111000100110",
"01010000010111001101100000111001",
"00101110100101000110000000110101",
"01111001100101110100111100111101",
"00000101010110001001000000001101",
"10111111101100101111111110011011",
"10111111001101110001000000100011",
"01010110010101011000010111000100",
"00101000100110010111011011000010",
"00101101011101010110000010100101",
"01010001100001011000101010001010",
"10111100111110010100111111100000",
"11000010000000110110111100000111",
"10100000101000100101110001011111",
"11011110010010011101001001110100",
"01101011100000101000010101000100",
"00010011011110110000111001100100",
"11010010000001000110111011111011",
"10101100111101110110111000001000",
"00111010100110000110100100101100",
"01000100010101101111111101110011",
"01011010111010001000100001101110",
"00100100000011001110101011101101",
"00001100001110010010000011111001",
"01110010101100010000000001001000",
"11001101111100010000001000000101",
"10110001000001111111011001011101",
"10010010011101001000111111010001",
"11101100100001011111110010010001",
"00011000110010011011111100110010",
"01100110001000100110101111011111",
"00001110010100011111000001100000",
"01110000100111000001010101011110",
"11111110000011100010101101011000",
"10000000111001100111110001011010",
"11000010101111001110100110010000",
"10111100001011010111010011000011",
"11100000101010011101001100000111",
"10011110010000001111001111001100",
"00010010010110011111111001101011",
"01101100100101100101000011110010",
"10011111100110011110001000001001",
"11011111010101001111000011101010",
"00111001011000001011011011111111",
"01000101100100011101001000000100",
"00110111110011110101000111111100",
"01000111000111100000111000010100",
"00000110001001001000011110011101",
"01111000110001110010100101011100",
"11010001100100100110010001001011",
"10101101010111111101011001110101",
"11000010111001101101011010110110",
"10111100000011011111001110110001",
"11010100111101001110010101100001",
"10101010000001011100110111000001",
"01110110100001011111101000001010",
"00001000011101001001010001101111",
"11010100010100111110001001101000",
"10101010100110101010011001111110",
"10110011010100101110010001101011",
"11001011100110110110000010111111",
"00010111110100001001110010011001",
"01100111000111010001001110010110",
"11010110010001000011100100000111",
"10101000101001101111111001101111",
"11001001100011100001010001101001",
"10110101011001101010000110001110",
"01010011100111111111001011100100",
"00101011010011001101110110010110",
"10110010000100111001000111101100",
"11001100110111100000110011110000",
"00111000010101110001101100011100",
"01000110100110000101010110010011",
"00110101010011010011111110011011",
"01001001100111111010011010000001",
"10010001111010011011001001011110",
"11101101000011000011011101000101",
"10010110100110110000111001100000",
"11101000010100110101010001110100",
"11110110111100000101001010001111",
"10001000000010000101100110100001",
"11011000110010110010101011000100",
"10100110001000010100100100110111",
"10010100101010000101111101100100",
"11101010010000101001110110110000",
"00001000111101110010000011110100",
"01110110000001001001100001001001",
"11010000101001011111011110001100",
"10101110010001010110111111010110",
"10010100001010001110001101001001",
"11101010110000100000010110110011",
"01001010011010001010010011111000",
"00110100100011001101100110100011",
"11000101100111011011000011000011",
"10111001010011111100110010101011",
"11000001110110000100011111010011",
"10111101000101111000000111000101",
"10111001101011100000000010010110",
"11000101001111000101000111000010",
"10111001011000111010110010011101",
"11000101100011111110110011000111",
"01111011011100100010110000000111",
"00000011100001110100111100001101",
"00111101011011110000011001111001",
"01000001100010010001011100010001",
"11100011011100101001100111010110",
"10011011100001110001000111001111",
"00011101110110111111110100111001",
"01100001000101001111001111101011",
"11100111011001101111001011010011",
"10010111100011011110001001101010",
"11100010001110110001101011100001",
"10011100101011110010000110110001",
"11001110101000110111100100001110",
"10110000010010000111001011111100",
"11101101111100100010110110111101",
"10010001000001110100111000011001",
"10000010000100011101001110110100",
"11111100111000001011010001100101",
"10110100111001011001110101100000",
"11001010000011101011010101100111",
"01000010100100010000000101000000",
"00111100011000011111101010000101",
"01000010001101000011011011100000",
"00111100101101011101001111110010",
"10011111111110110010000001010111",
"11011111000000100111101111110000",
"10010111010110100111011100110001",
"11100111100101011111110111011000",
"00011001100001001011100101101011",
"01100101011101101110001101000011",
"01000101011010101011001101110000",
"00111001100010111001110110110001",
"11000010011110001110101110001000",
"10111100100000111010010000000011",
"01000101101101100101000100010100",
"00111001001100111011101100101111",
"11010010001100100111001011000001",
"10101100101101111010000010100001",
"00011111111110010010110110010100",
"01011111000000111000000100011110",
"11111000010111101001111000010110",
"10000110100100110011000110110101",
"11111001110010111000001100101011",
"10000101001000010000001100101000",
"01111001000101111100001010111011",
"00000101110101111110101100111111",
"10011110100111001011000100101000",
"11100000010100010001111110100101",
"00100110010101011101011000110001",
"01011000100110010011110100001010",
"00010001011001000100110101101100",
"01101101100011111000011101100111",
"01010010110100001001000011100000",
"00101100000111010001110001101011",
"11110001000101011000100101110110",
"10001101110110110010000100111001",
"11010111101001010000001100000000",
"10100111010001101001010001110000",
"11001100011101001101001000100100",
"10110010100001011101100001000101",
"11011001001011100010010001110101",
"10100101101111000010101011110111",
"00000110001000001010000111011101",
"01111000110010111111111001101110",
"10010100101110010011111101111110",
"11101010001100001110001100011111",
"11000001100100101001010101011100",
"10111101010111111000101110001000",
"10101111011010010100000100111110",
"11001111100011000111101101000110",
"10100000100001010001011111010011",
"11011110011101100011010000100011",
"11100011110000000000101101100110",
"10011011001010101010000010001001",
"11101110110010011111011001111010",
"10010000001000100011111101101001",
"00000010000011100100101111100111",
"01111100111001100100011110011101",
"11011000000000010110010010010000",
"10100110111111010011111010001101",
"11100000111010001111011000101010",
"10011110000011001010100010001100",
"00010001010010101111100110001011",
"01101101101000010111000001010100",
"10111100111111100011011001001001",
"11000010000000001110011001111000",
"10100110100001010011100001000001",
"11011000011101011111100000110100",
"10001010110100001000001110101000",
"11110100000111010010011001100000",
"10000101110011001111010110110100",
"11111001000111111110000000010010",
"10000100110110011000111111111010",
"11111010000101101001110101000000",
"01010111110001001000101010000010",
"00100111001001101011100100110100",
"00100010110001000001000001101001",
"01011100001001110010000100000111",
"10101110111101011010101100010110",
"11010000000001010110001000010011",
"00111011010101000011010010001011",
"01000011100110100110101010100010",
"01100011010110111110100111110001",
"00011011100101010000000011111010",
"10101011001001100100100100110010",
"11010011110001010000111011100101",
"01100101110001101010001010001011",
"00011001001001001111011101001000",
"00100100110000110000000001111110",
"01011010001010000000101000010100",
"00111111110010001100011001100110",
"00111111001000110011010100100100",
"11111001011100100001111100010111",
"10000101100001110101011001001000",
"11110110011001000111000000010001",
"10001000100011110111000110100011",
"01011001010010000000100100001100",
"00100101101000111100111110100001",
"11101000010000010100101011011101",
"10010110101010011000011010001000",
"00001000000111101111110101010111",
"01110110110011100001100111111101",
"01110111101101000110100010000000",
"00000111001101011010000111101110",
"00101001000111110101000001110000",
"01010101110011011010111001111101",
"11100111000100010101001110011011",
"10010111111000010111101001110110",
"10011001001101101000001111000100",
"11100101101100111000100101000101",
"11010010011001110111110010101001",
"10101100100011011000110111101110",
"00110011110001101010000001000001",
"01001011001001001111100100101111",
"10010001111011010011100011000010",
"11101101000010100010000111100100",
"11110001001000001011010100011011",
"10001101110010111110011000000001",
"01101010111111000010100011001111",
"00010100000000011111001100010101",
"11101110110001010111011101100100",
"10010000001001011111000100110011",
"11110111101001001110110001100010",
"10000111010001101010111110101100",
"10010001000100101110110111011100",
"11101101110111110000010011100010",
"01101100011110100011100100111011",
"00010010100000101111010001110100",
"01101010001110101100001000111001",
"00010100101011110111010011010101",
"11001000011111001000111111101111",
"10110110100000011011111000000110",
"10111100101000101000011100010000",
"11000010010010011001110101110001",
"11010010001111010100011101101011",
"10101100101011010001111011000000",
"00111000011000111110001010101000",
"01000110100011111100101010100101",
"00110001101001010011100001011010",
"01001101010001100101010001010000",
"11001111010101011001100110110111",
"10101111100110010110100001101101",
"00100110001001010001111010111100",
"01011000110001100111001100010101",
"00111001110100000001101110011101",
"01000101000111010111010011110001",
"11100010000010010010001101101011",
"10011100111011101111000011110001",
"00101111110001100011001011001011",
"01001111001001010101010001001100",
"11000000110101001000011001010011",
"10111110000110100010111100110111",
"11110111110010100011101101101111",
"10000111001000100000100000010111",
"10000110110000110100000010101011",
"11111000001001111101001011011001",
"00100110100000101100111100101000",
"01011000011110101000000010010011",
"01110011001110000010000000110011",
"00001011101100011111011100011110",
"11000111111110001111110111111110",
"10110111000000111001101001000000",
"00000011000101110101000011110011",
"01111011110110001000110110011011",
"01111011111001011010100010010010",
"00000011000011101010111001110010",
"01101010010111010101110010001111",
"00010100100101000000011110000001",
"00001110101000110011001101100100",
"01110000010010001100100010001101",
"10000101111000111111000110100111",
"11111001000011111100000100110000",
"10100000000011110100100111101101",
"11011110111001001010111101011111",
"11100001000101010000011100010011",
"10011101110110111110000011110001",
"01100100000110110110011111100001",
"00011010110100101101101010111101",
"00000100110100000011011001000100",
"01111010000111010110000011001010",
"10010000001000110111011010111000",
"11101110110010000111010111011010",
"10110010011011010100010011011100",
"11001100100010100001101011011000",
"11111110000111100010111101001100",
"10000000110011110010011001110010",
"00010000110010101101101101110010",
"01101110001000011000100001001000",
"10101100011011011111111101101101",
"11010010100010011010111010010110",
"10110101010111101000111111010110",
"11001001100100110011101100100001",
"10111111101101111010101111001000",
"10111111001100100110011111101011",
"11111001000000101000001001111001",
"10000101111110110001001111000100",
"10001101110010100111100100100111",
"11110001001000011101011010110011",
"11101111111001101101111110010101",
"10001111000011011110111000111101",
"01111010011001100111100110100110",
"00000100100011100010110100000011",
"10100001110100111110000110011111",
"11011101000110101010011100010001",
"01111001010100010010001101101011",
"00000101100111001010111001010100",
"10011110100110011010101100110111",
"11100000010101010011110011100001",
"10011001110100001110010000101101",
"11100101000111001101110111000100",
"11000011110001100001011001000110",
"10111011001001010110110000011001",
"00110110101010101101010000010110",
"01001000001111111101000101110011",
"00000101011011101010111010010000",
"01111001100010010100100110001111",
"11100110100001010100010000000111",
"10011000011101011110001001111001",
"11001011011110001010101100101110",
"10110011100000111100011000010100",
"00100110010000111010101101101000",
"01011000101001110111011101001101",
"11010100010110011011010010100111",
"10101010100101101000001111100000",
"01000110110011011010101101010001",
"00111000000111110101001011100101",
"10000010101001100000110011101010",
"11111100010001010101011001101110",
"00101100011111110101110000100011",
"01010010100000000101001000100011",
"10100001011110100011111010111110",
"11011101100000101111000110010010",
"11010100011100111101010010111010",
"10101010100001100110001101100000",
"11010100010000101000011101000011",
"10101010101010000111001011001101",
"00011000111011001011101111011001",
"01100110000010100110101011000110",
"10100001110010101010000111100001",
"11011101001000011011011000101011",
"10111010010100011001010001111001",
"11000100100111000101100111001111",
"10011110100101110001011110110010",
"11100000010110001101111110101010",
"10011111111010110010010110000000",
"11011111000010110101100111111000",
"01110001100111001111000100000110",
"00001101010100001100101010001011",
"00100001000000000010111110010110",
"01011101111111111010000011110111",
"11110110100101000010011110100100",
"10001000010111010010110010001011",
"00110111001001101100101001010000",
"01000111110001000111011001011000",
"01010111011111100001001000001100",
"00100111100000001111100011011010",
"01110100000101100101110111011101",
"00001010110110011110101110110000",
"00111011110101010101100000011000",
"01000011000110011001011110011101",
"01001111000010000100000001100110",
"00101111111100000111111100010000",
"01101110111010001111011111000011",
"00010000000011001010011110010101",
"11111000000110101111100011111111",
"10000110110100110111000110011011",
"00010110100010011001010100010010",
"01101000011011100010101110010000",
"10110001001111101110101001110111",
"11001101101010111010001011000100",
"11101101101110101000011011111000",
"10010001001011111010110010010001",
"00010000110010011010110011101010",
"01101110001000100111101010011000",
"00101011010100001100000111111010",
"01010011100111001111011101110110",
"10010001011011011111101001100011",
"11101101100010011011000110000000",
"10011100000110001010001100011000",
"11100010110101101010110111011101",
"10110100110011100100111101101111",
"11001010000111101101010000100111",
"10100111110010000000111000110111",
"11010111001000111100101101100110",
"11010000000011101001110110110011",
"10101110111001011100001110001010",
"00100101110000011111000011111010",
"01011001001010001111010101010101",
"01010101010101100000110010101001",
"00101001100110010001011000001100",
"11100100101110101011010110010000",
"10011010001011111000000010111010",
"00111110111001101101111111101000",
"01000000000011011110111000001010",
"11000111110110100110001000110000",
"10110111000101100000110001000101",
"00010110110011110010110001011011",
"01101000000111100010101011001001",
"01001000000010011000110111000000",
"00110110111011100011100000111100",
"00010110101110000010111000110101",
"01101000001100011110100110010101",
"10110011100111101001010111000011",
"11001011010011101010000010011010",
"01000010000101011011001101100010",
"00111100110110101110001111011100",
"11011000001101101010110110001010",
"10100110101100110110000000110111",
"01111011110111010000101010111111",
"00000011000101000011111001001011",
"00000101111100011101011110111110",
"01111001000001110111111000110110",
"10000110111111000001101101011111",
"11111000000000011111101000000010",
"00011100101000000111001111101110",
"01100010010011000011100011010100",
"00101101000000000000011000111000",
"01010001111111111111001110010001",
"10011011001011111011010010100010",
"11100011101110100111111001101000",
"10100011111110011010110111111010",
"11011011000000110011110101111110",
"00100110101101000101111111110001",
"01011000001101011010101010001100",
"11010011100011100001011110000111",
"10101011011001101001110001111111",
"00011001111000100110011011001001",
"01100101000100001011101111101001",
"11001100111100101011100101100011",
"10110010000001110000000001000000",
"00110010011010110101101010110100",
"01001100100010110011101001110111",
"00010111101100000000100101000001",
"01100111001110100010010011000010",
"10001011001011001100001010110111",
"11110011101111011010110001000001",
"11000100111110010100100000110110",
"10111010000000110111001100010001",
"10101101010010010110101001101000",
"11010001101000101011000000111110",
"11010111101100101100000011100100",
"10100111001101110101000001011101",
"11110001100000011010110100100011",
"10001101011111001011000011010010",
"11100000111101010010100000011100",
"10011110000001011010100101010110",
"10110101101110011001010101010110",
"11001001001100001001000101001100",
"01010000100001001000010111111001",
"00101110011101110100001100011010",
"10010000010010110100000100110110",
"11101110101000010011011101100111",
"11010000110100111011010000101011",
"10101110000110101100100001000101",
"01010111010111101100000111010101",
"00100111100100110001101000010110",
"10100101100011100110001101001000",
"11011001011001100010000111001110",
"10001110101111110000111110010100",
"11110000001010111000000101101101",
"11010011001011010001110100101000",
"10101011101111010100100100101010",
"01010110001011000000010001000011",
"00101000101111100111111001000010",
"10100111001101000101101011000001",
"11010111101101011010111111000110",
"11000100101000101110001100001101",
"10111010010010010010101110010101",
"01000100101111000011011100111100",
"00111010001011100001100100011011",
"00101101000000111111010111101100",
"01010001111110000101000100000101",
"10100101001001111000111110011101",
"11011001110000111000111100000011",
"11111011000111011101010001100100",
"10000011110011111001110111000010",
"00101100101001111100010000100001",
"01010010010000110101000111001100",
"00010100000100011110011000001110",
"01101010111000001001100000100010",
"10000001110000001011001110110010",
"11111101001010100000101110000101",
"01110001101010100111111000001110",
"00001101010000000011001000111101",
"11011011010111001100100001101100",
"10100011100101000110101011010100",
"11110110111101100011001110010000",
"10001000000001010001100000100011",
"10111010010010100110100010000010",
"11000100101000011110010000000001",
"11110011011011000100100001100000",
"10001011100010101010111001101011",
"01000110110111111010110101101110",
"00111000000100100111111100100101",
"11111000010101001010110000010101",
"10000110100110100001001111010111",
"00101010111100010001001110011111",
"01010100000001111110110001110000",
"11011010010000011010101100100110",
"10100100101010010011001001000000",
"00101110111000111101110010011000",
"01010000000011111100111001111001",
"10001100000111000100001011111100",
"11110010110100011011001100010110",
"00100101110010110100010000100001",
"01011001001000010011010100010111",
"01011010001010000010001111101111",
"00100100110000101110001010000010",
"10111000000100011000000100011010",
"11000110111000010011001111110101",
"01001111100111110101001001011101",
"00101111010011011010110000000000",
"10010010100101110011000101000010",
"11101100010110001011101011111111",
"10001100011001101001110010101010",
"11110010100011100001011101101100",
"10001010010100110001000001001110",
"11110100100110110100000001110000",
"11101110110111110010010101100100",
"10010000000100101101100001110100",
"00001001000100100001001101100000",
"01110101111000000101001001110011",
"01010010000101001111111001111100",
"00101100110110111110110110011111",
"10101011111000111011101001101000",
"11010011000011111110010000010000",
"10111110000001011100100011111101",
"11000000111101001110111000011011",
"10000111011000010011100110110011",
"11110111100100010111110101100101",
"01000110100000100001100011100011",
"00111000011110111101111110001001",
"10011111100011010001010100110101",
"11011111011010000100001010111110",
"00001010010100001000001010000001",
"01110100100111010010011100111111",
"01011001110110000111001100111111",
"00100101000101110110001101100000",
"10010111110010110110000110011001",
"11100111001000010001110110111011",
"01010010101100101011000001101110",
"00101100001101110110000101000000",
"01001011101111000010100100100101",
"00110011001011100010011000100100",
"00101000101101001000010001100001",
"01010110001101011000010111100001",
"11010011001111011101101101011111",
"10101011101011001001011111010111",
"11011011011111111001011000001011",
"10100011100000000011010100010000",
"11110111101001010000110110000000",
"10000111010001101000011111001110",
"00100100011010000110111010001000",
"01011010100011001111101010100000",
"00110100100000110110101000111001",
"01001010011110010101100011111101",
"00010100001000111011011010001101",
"01101010110010000010011110110001",
"10100111001000001111011011111000",
"11010111110010111001001010010011",
"10001010110100001010011101011001",
"11110100000111010000101101111111",
"01010001110010100000011010001101",
"00101101001000100011001010000001",
"01000000010000010110101110111010",
"00111110101010010110100110111011",
"11101111101101100001010111100100",
"10001111001100111111010110011100",
"11000000100100110010111101111111",
"10111110010111101010000101101110",
"10101100000000111101001101010010",
"11010010111110001001001000110011",
"11101110111011000010101101110011",
"10010000000010101011111101101000",
"01111000100011111100000110011101",
"00000110011000111111000011111010",
"11001111111000101100001001000111",
"10101111000100001000000110000011",
"01001010101010000100010010000100",
"00110100010000101011110011000101",
"00001101111010101001110111000000",
"01110001000010111010101010011001",
"00001111111101000000000110111101",
"01101111000001100100101010010110",
"00001100000001110101111000000001",
"01110010111100100001000101001000",
"00000010100111110011010100111001",
"01111100010011011101000110100101",
"10110111000000001001111100101100",
"11000111111111101100001100110010",
"10111011101100000000010011001111",
"11000011001110100010100101110110",
"00010111011000110011110000001100",
"01100111100100000011010000010011",
"01101100001011110000001100010011",
"00010010101110110011101110011101",
"01101001100101001001010001101011",
"00010101010111001000101010011111",
"01110001101111101000011010111111",
"00001101001010111111110010011001",
"11100011011001101001000001110101",
"10011011100011100001111011110010",
"10111101011011011010001111010111",
"11000001100010011110001110100110",
"00010101100000100101011010001000",
"01101001011110110110100001101001",
"01101001111100110110101110111101",
"00010101000001101001110101010110",
"10000001110010110000001001110001",
"11111101001000010110100101000000",
"00010000110001110111000100100010",
"01101110001001000100110001100111",
"01110110111010010000001001000110",
"00001000000011001010000100111101",
"11000010000010001010110001111010",
"10111100111011111100000011100010",
"11100101001100101101111011010110",
"10011001101101110011000110101100",
"10100011000110110111010011010101",
"11011011110100101100100100101100",
"11101110011010000000110111100100",
"10010000100011010011010101010111",
"01011110000001001100010010001000",
"00100000111101101100111010011001",
"01101100010001011000010100000001",
"00010010101001011110010111000011",
"01011101011011111111000110110110",
"00100001100010001001000010101010",
"10100110000110001110000010010100",
"11011000110101100101011110000110",
"11101100111100001101001010000110",
"10010010000010000001000100101110",
"11011011110100100010110011110010",
"10100011000110111110100001100010",
"01110011011011001110011010100010",
"00001011100010100101000111000111",
"11100111110110000100000111011111",
"10010111000101111000010111110001",
"11111010011000010100100011110001",
"10000100100100010111001110001101",
"10000100111011011000100101000101",
"11111010000010011111001100010010",
"00011001010110110010010111100001",
"01100101100101011000011001001001",
"01110100001110101010101101111110",
"00001010101011111000101000110010",
"00001011100111100001011101110011",
"01110011010011110100010110110010",
"00011010110000011000001010111011",
"01100100001010010101010110010111",
"11110110001000011001100111111001",
"10001000110010101100010100111100",
"11000010111110100000111011011111",
"10111100000000110000101010100011",
"10111000010000010011100001100111",
"11000110101010011001011010111011",
"10101100011011111101100101110100",
"11010010100010001001111001111010",
"11110010100100100110000001111101",
"10001100010111111101110001000110",
"11110101101100101001011011101011",
"10001001001101110111101101110010",
"10011011110100111101010100001010",
"11100011000110101011000001000001",
"10010100001010100010011000011111",
"11101010110000001001010110010001",
"11011110010101110110011010100000",
"10100000100110000010000000101011",
"01111100010010111100100111101010",
"00000010101000001100101101000010",
"10101010001110110010010110100110",
"11010100101011110001011110011110",
"10010100001101001111010010000100",
"11101010101101010001010101100100",
"10001011011001101000011000011011",
"11110011100011100010010101010100",
"00101111110111110110001001110001",
"01001111000100101011000001010010",
"00100111101111001011111010000010",
"01010111001011011001110001010100",
"01100011111011110011111100001110",
"00011011000010001111011010100101",
"10001100111100100011001010111001",
"11110010000001110100101101010000",
"11010011110010011011110011010101",
"10101011001000100110110111000110",
"01010100011100111000110100110011",
"00101010100001101000101011011000",
"01010010110000101011100000101000",
"00101100001010000100100010000001",
"00010100110000001010101011000010",
"01101010001010100001001101101000",
"10110011010001011010000110101011",
"11001011101001011100110110110011",
"11110010010000101010010000011011",
"10001100101010000101100111010111",
"00110111011101100011111111110010",
"01000111100001010001000101110001",
"11110100111000011111100000110001",
"10001010000100010000001010111111",
"10000100001101010101110111010010",
"11111010101101001010110001000000",
"00101011010111000110000000000010",
"01010011100101001011000100100110",
"11010100111101100101101011110001",
"10101010000001010000001011011100",
"01000111011000001100100110010101",
"00110111100100011100010111110101",
"10111000010010110000011000110001",
"11000110101000010110011001000101",
"10110100100001101000111100011100",
"11001010011100111000010101111010",
"11011001110101000101010101111001",
"10100101000110100101001010110000",
"10111000011010101011110010110101",
"11000110100010111001100000101101",
"01111010110110101100111000000011",
"00000100000101011100001001010100",
"11110011111110100010111110100001",
"10001011000000101111100101111011",
"11010111000001000110111000000110",
"10100111111101110110111111010010",
"10111100001101000001001101011110",
"11000010101101011111011111001101",
"10110001101001011010101101000101",
"11001101010001011100101010111110",
"10011011111001110001011111111100",
"11100011000011011100101110011001",
"00011101000001010010010101111111",
"01100001111101100001101011011011",
"10100000011001111110010101110010",
"11011110100011010100110111111000",
"00101111111001100010111000000101",
"01001111000011100101101110111010",
"00111001101001001101010110100111",
"01000101010001101100101100010010",
"00000010100001110010101110010001",
"01111100011100100110101110011011",
"00001001101100100100011001011001",
"01110101001101111100111001011110",
"11110000001000110010011101010100",
"10001110110010001101011101100101",
"11010111000011000111011100000010",
"10100111111010010100100001010011",
"01110111100101011000111100011100",
"00000111010110110001100011110010",
"00011100010101010111110110011111",
"01100010100110010111110010011101",
"11001000001010011110101101111001",
"10110110110000001101100000001010",
"11110100010010101001100100100001",
"10001010101000011011110100100111",
"01111101101000111111101101010110",
"00000001010001111101001110111011",
"00110010110101001011011001010001",
"01001100000110100000110001101101",
"00001111000011000010111110011110",
"01101111111010011011111100100000",
"00101010010101000010001110000000",
"01010100100110100111011100001010",
"01110001000101000101111100100010",
"00001101110111001101100111010011",
"11111011001110000101101010000101",
"10000011101100011011111011010001",
"01011111000101101101101001111100",
"00011111110110010011011110101010",
"10101011101111101101010000000110",
"11010011001010111011011011110011",
"00111000100100011011011111011001",
"01000110011000001101111101011010",
"10100111000000011111011001001011",
"11010111111111000010001010010101",
"01100101110110010111100000100111",
"00011001000101101010110111000000",
"00011111000101010110001010010010",
"01011111110110110101101001000101",
"10100001001111111111001011100100",
"11011101101010101011011001010011",
"11001000111111101100011000000010",
"10110110000000001001110111000000",
"10101110110001001100101111010110",
"11010000001001101000000111011011",
"01101101110001111101110100110101",
"00010001001000111111001110010000",
"01100011001110011010001110001010",
"00011011101100001000001111001010",
"01000101111100111101101001111110",
"00111001000001100110000000110011",
"11110000011101100110111101010110",
"10001110100001001111011111011010",
"00100001101110011110100000111000",
"01011101001100000100001010010100",
"11001010100000100100111110000101",
"10110100011110110111010111110000",
"10001100010001000000001101000010",
"11110010101001110010110000111110",
"00011010101100011100100011010100",
"01100100001110000101000000100100",
"10010010011000100100101011010111",
"11101100100100001100110111001000",
"01010011111001001101001010100010",
"00101011000011110011001111011001",
"11100010111000011010111110001000",
"10011100000100010011000101101110",
"01100000000101111100111010111000",
"00011110110101111101101000110010",
"00010111001011010101001000001101",
"01100111101111010000111101100101",
"10111101011000011111001001001011",
"11000001100100010000011010001000",
"11101010110000011001111111111001",
"10010100001010010011110000000100",
"00011101011101010111011100110011",
"01100001100001010111111001000101",
"10011000100011111000010101001101",
"11100110011001000101000011000100",
"11111001001001100001000010110100",
"10000101110001010101000111101110",
"11110010111101001110110111100101",
"10001100000001011100100100011010",
"11001110110010110101110111001010",
"10110000001000010010000011000000",
"11001011001001110100111010000011",
"10110011110000111101101100011100",
"10110001101000010001100011011011",
"11001101010010110110011111000001",
"11000010111001101101011101010001",
"10111100000011011111001101010010",
"00001111011011100010100100001101",
"01101111100010011001011010000101",
"10011111100101100110001001011100",
"11011111010110011110010100101100",
"00001110101011010110001101001010",
"01110000001111001111110010011001",
"00011101000100010100011001111001",
"01100001111000011000111011011000",
"00000100011011110010001111111110",
"01111010100010010000011000100101",
"11110000000111001111001110011110",
"10001110110100001100011100010111",
"10010100011010101011000010010110",
"11101010100010111001111101100011",
"10101101111101111101010001101010",
"11010001000001000011100001000101",
"10110011011010000001000011000110",
"11001011100011010011001110010110",
"00110010100011110100001010000110",
"01001100011001001011101100110000",
"10100101000010101011100110000010",
"11011001111011000011010101111101",
"10010110001010101010000110000101",
"11101000110000000000101001001011",
"10111010001100110000011010001000",
"11000100101101110000100100001110",
"10001101001000111100010010011100",
"11110001110010000001011010000010",
"10111000101111010100000111001110",
"11000110001011010010001111100011",
"00111000001001110000000100010010",
"01000110110001000011010111101110",
"00100101010100111011111000010101",
"01011001100110101100000100000110",
"10101011011111100110011010001011",
"11010011100000001100111000000100",
"01011010001101010111010101010010",
"00100100101101001001010011011010",
"00100010110001100101001101100001",
"01011100001001010011100100100001",
"11111100110011100100010110001011",
"10000010000111101101101111000101",
"10100000011101011010111110011001",
"11011110100001010101111110100000",
"11101101110000011101101010010111",
"10010001001010010000100011011000",
"11000011000110010001110111101010",
"10111011110101100000000110101001",
"00010100111101001101110110111010",
"01101010000001011101000111110000",
"11001101101110000000110011010111",
"10110001001100100000100111010110",
"10011011001011001001000011011011",
"11100011101111011110001100001111",
"10101101110101011010111010001010",
"11010001000110010101100101111010",
"01000101001101001001111001100110",
"00111001101101010110101110111011",
"01000001001100111011011011000111",
"00111101101101100101010110001101",
"10001011000001000000111100010100",
"11110011111110000010000110111000",
"11000110000111010100101100010000",
"10111000110100000101001100000110",
"01010001000110000001101101001000",
"00101101110101110110110110001100",
"01100100010110001110111010001001",
"00011010100101110000110101010110",
"00111010001010110101111010100000",
"01000100101111110011011001100001",
"10001001111100100010100111101011",
"11110101000001110101000000111011",
"00011010000000101000100011101010",
"01100100111110110000011101100000",
"11001000001100101001101001001100",
"10110110101101110111011111111001",
"01111000110101010101110110001000",
"00000110000110011001001110110011",
"00101000111011100100111011011110",
"01010110000010011000000010110000",
"10000000111101000001100010100110",
"11111110000001100011110111111011",
"11000111110010011101001001111111",
"10110111001000100101110001010110",
"11011010100010010000101000010010",
"10100100011011110001110100100100",
"01110001100000000100000011100101",
"00001101011111110111111001111000",
"00110000100110001111010000110000",
"01001110010101100011110000001011",
"00011101101011111000100010101101",
"01100001001110101010110100011100",
"10101100000011101010111110000101",
"11010010111001011010011011011000",
"11101011111101001101000001101101",
"10010011000001011101100100110101",
"01010101011010001000010101011001",
"00101001100011001110110011001011",
"00101000011101000101101101101000",
"01010110100001100001100101001110",
"11010111011011010000000011100001",
"10100111100010100100001001110101",
"11000110100011011000100000100101",
"10111000011001111000011000011111",
"01011100110011100101111011010111",
"00100010000111101100100001001100",
"11111001001100111110110101001100",
"10000101101101100001111001001101",
"00011010000010111101101010101000",
"01100100111010100100110100100000",
"11100011011011011111011110100010",
"10011011100010011011001100011000",
"10011000110010001001011111011111",
"11100110001000110101101011111111",
"00110111001000001001110011010000",
"01000111110011000000010011011000",
"10100000110101110100101100101011",
"11011110000110000011001110010010",
"10010011000011110100101001101010",
"11101011111001001010111010011000",
"11011011010101001101010101100001",
"10100011100110011111010111110010",
"10001101000011010100001010011111",
"11110001111001111111100000010010",
"00010100100010111010011011010101",
"01101010011010101010010000010011",
"00000100100010100100111110110100",
"01111010011011001110101000101111",
"01001001010011111101001000000011",
"00110101100111011010110010110101",
"01111001100010000001000000101000",
"00000101011100001101010001010101",
"01011111011001010011000001101111",
"00011111100011101111100100111101",
"10010010001011000101110010101111",
"11101100101111100001110010001001",
"11001110110101011011101011000000",
"10110000000110010101000010110111",
"00010001110101110100101110100110",
"01101101000110000011001100111011",
"00101101100000101000011000100101",
"01010001011110110000110010110011",
"00000011111000011000100010110111",
"01111011000100010100101001101100",
"00100000011111010000110101101010",
"01011110100000010111110110110000",
"10111001100111001011111111110110",
"11000101010100010000101111100101",
"11100011101000110000001100111101",
"10011011010010010000001111011100",
"10010010110001001001011111110000",
"11101100001001101010110111010000",
"11111101011010101101110101111000",
"10000001100010111000010010110101",
"11000110010110110101110110000110",
"10111000100101010110000001011011",
"00011000110100111110110110011011",
"01100110000110101001111001010010",
"01111011111010101011000001111100",
"00000011000010111001111101110011",
"01110111111001000101100001010111",
"00000111000011111000000010001010",
"00000010111000001001001010000010",
"01111100000100011110100110110101",
"10110101100010000101100011110010",
"11001001011100000101001111000100",
"00010011011111010001100000001101",
"01101011100000010111100000111111",
"00100000011011010011100100101100",
"01011110100010100010000110100110",
"11101101001111111010100100011011",
"10010001101010101111100000001011",
"00011010100110011010011011111100",
"01100100010101010100001011000000",
"00010100001110101101110101010110",
"01101010101011110101101101011111",
"00101100001000110101011101011010",
"01010010110010001001110001011000",
"01111100011010110000110011111011",
"00000010100010110110100010000001",
"10011010100000111010011110101101",
"11100100011110001110010010011010",
"01001110101111100011001100110111",
"00110000001011000100100000100001",
"10101111000000010111111101111010",
"11001111111111010000100111101011",
"00101001111001010000100101110011",
"01010101000011110001000110010011",
"11011111111111110011110111110111",
"10011111000000000110000101001110",
"00101001111110010010110010110100",
"01010101000000111000000110010100",
"10011011010000100111101010010100",
"11100011101010000111110111001001",
"00101111001011010001111100010101",
"01001111101111010100011100001111",
"01000001111001101010111001101000",
"00111101000011100000110001111111",
"11010101001010001110011100111001",
"10101001110000100000000100101101",
"01100111111111101001101011010110",
"00010111000000001011001110010000",
"10110000010000111010011011100110",
"11001110101001110111101100101000",
"00110011100010011100001000100110",
"01001011011011011101110110100000",
"10111101101011101111011000111001",
"11000001001110110100100101011110",
"10010010010101100010000110001001",
"11101100100110010000011100011111",
"01101111011100110111010000011001",
"00001111100001101001100010110111",
"01001001010010011010100000100000",
"00110101101000100111111001110100",
"11000100110010000100111001011100",
"10111010001000111001011011110010",
"01010011010010110011100000001101",
"00101011101000010011111010101100",
"01000000001000001001010010110001",
"00111110110011000000111100101010",
"10010100011111010001000110111111",
"11101010100000010111101101111001",
"10001011001011100000110001010011",
"11110011101111000100010100001110",
"00010110111100111000000010011100",
"01101000000001101001000111001100",
"10000000100010100101111111011010",
"11111110011011001100111010001001",
"11111101000001010110001010001010",
"10000001111101011010101000111011",
"10111011001011100001011010011010",
"11000011101111000011100111110001",
"00011000000110111101011101100111",
"01100110110100100100001111011001",
"11100111100111000011111100110100",
"10010111010100011011100000101001",
"10101111111100000100000110111101",
"11001111000010000110001100101101",
"00101011010100101011001100001110",
"01010011100110111000010100100110",
"11011111011001010011100010100010",
"10011111100011101111010000011111",
"11101111001000000010110001111100",
"10001111110011001001001111101100",
"11011000111101111100111001110111",
"10100110000001000011101101110010",
"00100000111110100000100001011110",
"01011110000000110000111000001100",
"10100010100101011101001010101001",
"11011100010110101011011000101010",
"01011111100011010111110010001001",
"00011111011001111001100100011111",
"01001011001101000101111001110100",
"00110011101101011010110000001100",
"11100110110100100111000010111100",
"10011000000110111011011000101001",
"00100101000101101011010001000100",
"01011001110110010110111011000000",
"00111011000000100000111000010110",
"01000011111110111111010001110100",
"00111101000100000001011110101001",
"01000001111000110110100011011011",
"00000111001000000001010000101111",
"01110111110011001011001011111010",
"11100001101000011110001000110000",
"10011101010010100110101011001000",
"10100000110100011000100010011101",
"11011110000111000110001010101001",
"00010100000001111000100011010001",
"01101010111100011100010011010001",
"11010011110110001000011100110011",
"10101011000101110101010101101101",
"01100110111010100110001011010011",
"00011000000010111100110110110110",
"10011100000110111010001000110110",
"11100010110100101000101110110110",
"01110110111000010010111010001001",
"00001000000100011000010010011011",
"01101100001001010011011111001111",
"00010010110001100101010011110111",
"00011110001100000100011110100011",
"01100000101110011110001011100010",
"01010000100010011110010110011010",
"00101110011011011010000001111001",
"00110110011011100011110100110100",
"01001000100010011000101011100010",
"01001011100011001000010100101001",
"00110011011010010011000011010101",
"10011110101110010010011011101100",
"11100000001100001111101010011000",
"11111101101000010000100001000111",
"10000001010010110111110010110010",
"01111100101111101011011111101111",
"00000010001010111101000000111110",
"10110000111101010010110110100101",
"11001110000001011010011001010001",
"11110011011111010110111111011010",
"10001011100000010100101101100100",
"11101111111100101011111000001101",
"10001111000001101111110110101000",
"00011101111010101111000111101111",
"01100001000010110111100010001101",
"01111010111100011011101000011110",
"00000100000001111000111011010001",
"10000110110000111111100011110000",
"11111000001001110011010100001100",
"11000100101101111000011000001101",
"10111010001100101000110010011001",
"11010100001000110000011011101001",
"10101010110010001111111101010101",
"10010111000111000010100010101011",
"11100111110100011101011001101101",
"01111100100011110111001000110101",
"00000010011001000110111100101000",
"01011011101101111111010010100101",
"00100011001100100010000101000001",
"00011111000000100110010010011100",
"01011111111110110100110101000100",
"10001110100000101010000011100010",
"11110000011110101101100101010000",
"10101101110100110000110100001101",
"11010001000110110100001011010101",
"00011001100001001100101000011110",
"01100101011101101100010000110111",
"00010000111001001100010110100000",
"01101110000011110011101111111101",
"00001000111100100101111100011011",
"01110110000001110011001010001010",
"00011100010000001010111000000111",
"01100010101010100001000010000101",
"00001011111001110010111000100101",
"01110011000011011011111000000010",
"10111100101100000110001001101001",
"11000010001110011100011010101011",
"10111111000000001111010010111000",
"10111111111111100001101000110001",
"00011101111001100100010010011000",
"01100001000011100100110111000101",
"01000001000110011000001011010011",
"00111101110101010111010011111100",
"00110100100101010011100010100011",
"01001010010110111001011111101010",
"01100100010111001001101000001111",
"00011010100101001000101000000101",
"00111111110110111011100111000100",
"00111111000101010010000110100101",
"11100100001000100101101001000010",
"10011010110010011101010100010101",
"11100111010110010000100010000010",
"10010111100101101111101101000011",
"10011100100110011010100111101010",
"11100010010101010011111010101111",
"00111111101111011101101010001011",
"00111111001011001001100010011000",
"00000000100110000110101111001100",
"01111110010101101111101110111111",
"10010100000011111001111101101000",
"11101010111001000010011101000100",
"11000001100101010101011011001111",
"10111101010110110110101110001100",
"01010111000001001011100111001001",
"00100111111101101110001010010100",
"00100110110011111011010111010001",
"01011000000111011100001000011100",
"11000001101110100001010010010001",
"10111101001100000001100010010010",
"00011001101111100010100101001000",
"01100101001011000101000100100001",
"10110110101111110100010111101011",
"11001000001010110101000010110100",
"01011011000010010100001011100011",
"00100011111011101011101000101010",
"01011011001100000110111010101110",
"00100011101110011011100111000000",
"01111001110000110001101100001000",
"00000101001001111111001100111001",
"01010110001111110110001000101011",
"00101000101010110011011101101010",
"11010111101101011000110010111111",
"10100111001101000111110110001101",
"01001100011110110011100011111011",
"00110010100000100110111100100011",
"11100100101101010111000001101000",
"10011010001101001001100110111110",
"01100000001000111010000011110001",
"00011110110010000100001000100000",
"01101001111011001011111010011011",
"00010101000010100110100100101001",
"00011000101110111101110101011110",
"01100110001011100110110001100011",
"10011111111111101011000011111000",
"11011111000000001010100001100000",
"11010110111101110010011011100110",
"10101000000001001001010100011001",
"00000100010000011000110110011000",
"01111010101010010100110000010110",
"01100100100011000101110011101110",
"00011010011010010111001110101011",
"10111111000010001011001000011001",
"10111111111011111011011100000110",
"11010110000111001011001101111110",
"10101000110100010001110010000111",
"11011010011110101001110001111000",
"10100100100000101100000010011001",
"10100010000110110010010111100011",
"11011100110100110011010001101101",
"01110011110101101001100101011101",
"00001011000110001011000110101101",
"11101010100110100111110001110011",
"10010100010101000001110000010010",
"01001101011000101000111010000111",
"00110001100100001010001010000101",
"11100010111111111000110101100111",
"10011100000000000011100101100110",
"00000100001010010101101000110110",
"01111010110000010111110101110011",
"10101010110111010000111011000000",
"11010100000101000011101110011100",
"01100100110111000010011000011000",
"00011010000101001101100001000011",
"00101111000001111001000100110101",
"01001111111100011011010111011010",
"00000011001001000111111101001101",
"01111011110001110011001101101101",
"11100110100100111001110010011010",
"10011000010111011111110011100000",
"01110110101101000000100001001010",
"00001000001101100000001011111111",
"01000010011001101110000001101001",
"00111100100011011110110110111011",
"00001010101101011001100101011001",
"01110100001101000111000100000111",
"11110100001111010111100101000001",
"10001010101011001111000100111000",
"01001001110100001011011000010101",
"00110101000111010000000001101000",
"00111001011011011110110101010010",
"01000101100010011011100100010000",
"00001110101100110010011100110010",
"01110000001101101110011110101110",
"10001001001100110111010110001111",
"11110101101101101001011111010000",
"11011011000111100001111100110100",
"10100011110011110011101110001000",
"00001110001011011011010010101001",
"01110000101111001010010000010010",
"10101111010101100011000101001111",
"11001111100110001111101111011010",
"01001101010111011001001000111011",
"00110001100100111110001110100110",
"11111100101000111010111110000111",
"10000010010010000011000001000111",
"00011001000011010010111001111000",
"01100101111010000001100100101111",
"00000010011000111101101110001101",
"01111100100011111100111100100001",
"10000111001011100011101110111001",
"11110111101111000001000111010111",
"11001010110000001100010010011010",
"10110100001010011111110010011011",
"10101110110101001001111000111011",
"11010000000110100001110111100001",
"01100010000110001011000000001011",
"00011100110101101001101110101000",
"00111010101001101001001111000101",
"01000100010001001011011010101100",
"10111001011010101011011010100000",
"11000101100010111001101111001011",
"01101001100100001011010110010010",
"00010101011000100111000010110100",
"00011000000111001110101011011101",
"01100110110100001101001010111101",
"00100100001100111001001110001100",
"01011010101101100111100101010010",
"11011110111101110010111000011001",
"10100000000001001001000100111100",
"01010010100000101000001101111100",
"00101100011110110001000111010001",
"01101011011011000000101110011110",
"00010011100010101101001000011110",
"10100010011111111011011011010000",
"11011100100000000010010010100010",
"10011100010001010011100100101001",
"11100010101001100010010110001111",
"01100111110101111110100111111001",
"00010111000101111100001110100000",
"00111011001011011011000001011011",
"01000011101111001010100010111111",
"00010111110000001111100010001101",
"01100111001010011100111011011000",
"10111000100110110100000111010101",
"11000110010100110000111001101001",
"01011011011001001101001011101001",
"00100011100011110011001110101100",
"01101001101001111010111001000101",
"00010101010000110110101101000011",
"01000110100111010101100000000000",
"00111000010100000100000111100101",
"10001010000111111110011111000110",
"11110100110011001110101111010100",
"11101011001100000100001010111000",
"10010011101110011110100000010010",
"00100010111100100011100010110101",
"01011100000001110100011111111000",
"00010101011101111101110010110101",
"01101001100001000011001111011001",
"01000001110001010001111001111001",
"00111101001001100011110000001110",
"10010000001101101100011000110110",
"11101110101100110100100000000001",
"10000111110110100111010111101010",
"11110111000101011111111010111001",
"10010101010000001110010100111100",
"11101001101010011101111111011001",
"11101110010000110110001001010000",
"10010000101001111011010111110011",
"11000010110010001100001111001001",
"10111100001000110011011101000100",
"01101100000111101111010011101000",
"00010010110011100010010011101101",
"10101111010111111000011110100001",
"11001111100100101001011111101011",
"10100001000111110101001100011111",
"11011101110011011010101100000110",
"10111111011011100010100010011110",
"10111111100010011001011011000101",
"00100000110011111100000100111001",
"01011110000111011011100101110011",
"10101101110110010110011001001011",
"11010001000101101011101000100001",
"10110110001110011000111000110001",
"11001000101100001001100000011001",
"01001101001011000111101110100011",
"00110001101111011111101001101011",
"00101000011011010111111101001000",
"01010110100010011111100011011111",
"11011011000101010010110110110100",
"10100011110110111010100000000010",
"11001010100111101011100010001010",
"10110100010011100111001101010100",
"00010111011000111100011111011001",
"01100111100011111101101110010010",
"10011110000000100111000011110010",
"11100000111110110011010110000000",
"01110110100110001101110110000111",
"00001000010101100101101111001101",
"00101001101111010111110001001011",
"01010101001011001110111001110010",
"10110101101101101110010111101101",
"11001001001100110010100011101010",
"10010011111010110101110110100111",
"11101011000010110011100010111001",
"00111010100101101010011111110000",
"01000100010110011000000010001011",
"01101111110110101100100000011010",
"00001111000101011100011001100000",
"10111111110100011011001000101011",
"10111111000111000100001110101011",
"00111011100110100011001001010011",
"01000011010101001000001000001001",
"00000110101101001100000101111010",
"01111000001101010100100010000110",
"00001111011101011010011001000101",
"01101111100001010110010010110000",
"11101011011010110000011001001110",
"10010011100010110110110001110111",
"10011001010101001101111010000011",
"11100101100110011110111101010111",
"01010101110101101100011111100100",
"00101001000110001001000010011001",
"00001000100000101110110101001101",
"01110110011110100100011011100111",
"11011101010111010101001101110010",
"10100001100101000000110110011010",
"00111000011111010110110000100101",
"01000110100000010100110101001001",
"00011100111101110100000011110000",
"01100010000001001000011100100010",
"00011010111011000101111110010101",
"01100100000010101010000011001110",
"10000001011100110111101010010011",
"11111101100001101001010100100010",
"01010001100100101011100101101111",
"00101101010111110101010010010010",
"00011011011100011011000100000010",
"01100011100001111001001111101101",
"10101110111100000100010100110101",
"11010000000010000110000100110101",
"10000111111011001110100111111010",
"11110111000010100100111111010011",
"11011111110100101001000101001011",
"10011111000110111001111000010110",
"01100100110001110100011101110001",
"00011010001001000110111011000111",
"00000001111011010110010000111001",
"01111101000010100000100010011001",
"10000001010001110101011001110011",
"11111101101001000110001001100110",
"00101110110101001100110001010001",
"01010000000110011111110010000000",
"11001011100111010110010011110100",
"10110011010100000011000011000001",
"00001000111001100000111010010101",
"01110110000011100110111100101110",
"10010011010011001110111110000000",
"11101011100111111110010011101001",
"00000001100100100110001100010010",
"01111101010111111101100001010011",
"10001101110011000100010010000111",
"11110001001000000110101010111110",
"00000111110100100001100101010000",
"01110111000110111111011011110100",
"10100111010001011110101001010110",
"11010111101001011001000011010011",
"11010000100001001110101111011001",
"10101110011101101000010110011000",
"00101011000001111101110101011011",
"01010011111100010010111001100001",
"00011001110000110111111010101110",
"01100101001001111001110110011101",
"00110101000110100011011110111101",
"01001001110101000111101010010100",
"01001010010101110101011110010101",
"00110100100110000010101011001011",
"01000100110100111010011110010100",
"00111010000110101101000101111010",
"10010111111111011010010100100010",
"11100111000000010011000000111011",
"10100100000010001110011111101100",
"11011010111011110101100011001000",
"01001111111001010100000111000111",
"00101111000011101110111001101100",
"11010011000001001001000100110110",
"10101011111101110010111000100100",
"00111011011000101011110111101100",
"01000011100100001000010001001010",
"10011010001011101100101100011000",
"11100100101110110111011110010100",
"10010110100101011011000100100110",
"11101000010110101110011100100000",
"11011001011100111110001110100110",
"10100101100001100101101100100111",
"10110111001110101100111010111010",
"11000111101011110110100100010110",
"11110111110011001001110100110110",
"10000111001000000010010100110110",
"01000011011100010110100101010110",
"00111011100001111011110000101101",
"00000111001101001110101110100001",
"01110111101101010001111001001001",
"01010101110010010100000111101000",
"00101001001000101101000011111011",
"11010110110010101111011111111110",
"10101000001000010111000110010000",
"01010110001100001010001010001100",
"00101000101110011000001100110111",
"01101100011001010101010101001100",
"00010010100011101110001001000001",
"01100001101110011001110110011001",
"00011101001100001000100101110000",
"10110101000000001011100100100010",
"11001001111111101000111111010001",
"00001010011010100010111110111110",
"01110100100010111110110000110100",
"01101110010101101100101100001111",
"00010000100110001000111001011001",
"11111000011011000110100100000011",
"10000110100010101001101101000110",
"01001100100101000000101001110101",
"00110010010111010101100000100101",
"10100011010101000100011010101100",
"11011011100110100101110101110010",
"11010010100110100001101010100111",
"10101100010101001010001010101110",
"10001011100011101001001111000010",
"11110011011001011101001110001111",
"10111101111101010101111001110101",
"11000001000001011000101110111011",
"11110011010000000110110000000001",
"10001011101010100100101011100000",
"01001111000100101010001011000001",
"00101111110111110111011100011100",
"10110011110111110011100111011010",
"11001011000100101100101011111111",
"01100101101010100000001110010010",
"00011001010000001011110010110101",
"00010011011100011000110011111100",
"01101011100001111010100000100101",
"00110000101100101100110001011110",
"01001110001101110100010010011001",
"01111001000000101000000010001101",
"00000101111110110001011101110110",
"11010000011101111001000001110110",
"10101110100001000101110010010000",
"11101100001111101001111001111011",
"10010010101010111110011100101111",
"00101000000001011010101100100001",
"01010110111101010010010011010001",
"01000011101110101101011110111011",
"00111011001011110110000010100010",
"10110110100010110101010000101000",
"11001000011010110010111101001111",
"11111000011010001000111011000110",
"10000110100011001110011100010101",
"00000010001100000000001001001010",
"01111100101110100010110000100000",
"10011111001100001111001011001100",
"11011111101110010010111100010100",
"00010110101110101010000111101100",
"01101000001011111001001100110010",
"11010011111001000000000100011100",
"10101011000011111011011101110001",
"11011100011111001100001011001110",
"10100010100000011010001111101001",
"00001011000100001000100111111011",
"01110011111000101011010011111110",
"10101000000001111100101000011101",
"11010110111100010101000010001110",
"00001001100010100110011110001100",
"01110101011011001100000101011110",
"11100110111101000101110100010101",
"10011000000001100001100001100011",
"10001001100000011110110011110010",
"11110101011111000011010010111001",
"10000101111110011001100001100100",
"11111001000000110100100011010111",
"11110110001110100100100100010001",
"10001000101011111110011011110001",
"01011010011010111001001011101100",
"00100100100010110001100100111101",
"00100010100110001111100100011100",
"01011100010101100011010100100111",
"00100001000001000011111100110011",
"01011101111101111100011101101110",
"00011010000111000101010111100100",
"01100100110100011001100110111010",
"00011110111110001010101001101010",
"01100000000000111100011001111011",
"01100011010110011010001000111101",
"00011011100101101001000010011100",
"01001011101111101010011101111110",
"00110011001010111101111100001111",
"00011011100000001001000100000100",
"01100011011111101101111100111111",
"10111111000000001101111001010001",
"10111111111111100100011001011101",
"01101010011000100011000010101101",
"00010100100100001101111010001000",
"11000101000100110011000111110110",
"10111001110111101001110110110011",
"10111111110000110011111011101010",
"10111111001001111101010001011011",
"11110110011110011000000001010011",
"10001000100000110101010110000001",
"11100011011100110111110010010110",
"10011011100001101001010000000110",
"10111111000001011011011101001010",
"10111111111101010000111010000110",
"00101010011100100101110000111101",
"01010100100001110011010000100011",
"10010011101000101110011001110011",
"11101011010010010010011101100010",
"10101010011010000011000101001011",
"11010100100011010001111111001111",
"11101000000011001101110100111011",
"10010110111010001001111100001001",
"11010111110110110110011100100101",
"10100111000101010101100111001110",
"01111101110100011100111111011111",
"00000001000111000010110110001100",
"00111100101110001101001111111100",
"01000010001100010100101000000010",
"01110010011100101010110010111100",
"00001100100001110000011101001010",
"11110001110010111110000110101010",
"10001101001000001011100010000111",
"10011000011111000011001101111100",
"11100110100000011110110110010101",
"01010000000110101010101010010001",
"00101110110100111101110011010100",
"01101111111001010100000100000000",
"00001111000011101110111011101000",
"00100001100001001001111001000011",
"01011101011101110001010111010001",
"01000011000001110100001110011011",
"00111011111100100100000010000110",
"00101101000001101000001100111110",
"01010001111100111001101011110110",
"11111001111110111001111111000100",
"10000101000000100011100111011100",
"10111010100001001111010100110001",
"11000100011101100111010001000101",
"01110101010100001000111101011000",
"00001001100111010001110110010010",
"11101000111010000101100000111110",
"10010110000011010000100000100111",
"00101001100101110101101000010010",
"01010101010110001000000010001110",
"00001000011000001111111111100000",
"01110110100100011010001011001000",
"00110000010010101001111101111100",
"01001110101000011011100000010101",
"00111110100010011001001100001110",
"01000000011011100010111100001101",
"10101100010001110011011110101010",
"11010010101001000111101111001101",
"01111110010001001001001101111110",
"00000000101001101011000110010101",
"10000001001100011100010100000010",
"11111101101110000101010000011010",
"00011101000000101101110110001100",
"01100001111110100110010100001000",
"00010100111100110110100011110011",
"01101010000001101001111011100001",
"01000100011011111100001110011000",
"00111010100010001010101011101110",
"00011111000100011101000101011110",
"01011111111000001011011111111111",
"01000101011101000100110001100111",
"00111001100001100010000110001011",
"00110010000111111011000010001000",
"01001100110011010011001010111000",
"00111101011100010100001000110010",
"01000001100001111101001000110010",
"00100010100010110001010000000101",
"01011100011010111001101111000100",
"11110100100111000011011001011110",
"10001010010100011100010000000110",
"00001101000100111100001010001110",
"01110001110111011100001111011011",
"00110010011100101001110000100101",
"01001100100001110001000010000110",
"11110111110100001110001011011010",
"10000111000111001101111011000010",
"01011111011101001110001100110001",
"00011111100001011100111011110011",
"10101110010100000100001001000000",
"11010000100111010101011110111011",
"01101000110110111000010110101010",
"00010110000101010100010100001011",
"10101100000110001011010010111110",
"11010010110101101001010100001101",
"10100000100110010000110101000100",
"11011110010101100001100011110001",
"01000100011001011101111100000111",
"00111010100011101000110010100101",
"10011001000001101100101000111111",
"11100101111100110001101010100011",
"01010110011111110001011110110011",
"00101000100000000111010010010000",
"11111100100001010010000110000111",
"10000010011101100010001000110010",
"11011110011101000101100000111111",
"10100000100001100001101100001010",
"00110000000011110000100000011011",
"01001110111001010001100010011100",
"11100000010011111111111000101010",
"10011110100111011000101100111101",
"01001101001000011101101001011011",
"00110001110010100111010010010011",
"00100001101010000111010010110111",
"01011101010000101000010100001101",
"00101010110000100010001011000011",
"01010100001010001100101000000001",
"01110000100100001010010110110011",
"00001110011000101000100110001100",
"10111101100100010111001000010110",
"11000001011000010100101100110101",
"11100111111100000111110010100011",
"10010111000010000100000111000110",
"11001110011000101110111100110101",
"10110000100100000110010011100111",
"10101100010010110101101011111000",
"11010010101000010010001011111100",
"11010101000101010100111100010010",
"10101001110110110111011011101011",
"11010100000001001100110101010101",
"10101010111101101011111000111110",
"01010100001010001110101001100100",
"00101010110000011111110110001010",
"11001100100101110010111111111000",
"10110010010110001011110011011000",
"10110011001000101010110101000011",
"11001011110010010110111000011001",
"10001010101001000110111110100101",
"11110100010001110100011001100100",
"10101100000010101111010001111011",
"11010010111010111101000100111110",
"00000111110111001111001111011000",
"01110111000101000100110110101001",
"01011000010110000010111010000111",
"00100110100101111001001101111111",
"01111000110000010100010101010110",
"00000110001010011000101101100001",
"11000010111111101100000000100010",
"10111100000000001010000010111000",
"00001101010100010101011100111110",
"01110001100111001000011110001010",
"10001000001100101101001011111100",
"11110110101101110011110111010000",
"10100110111111010010100111111001",
"11011000000000010110111100010101",
"10001001010010110000010101000010",
"11110101101000010110011100000011",
"01000101100100011011111010101010",
"00111001011000001101010011010101",
"11000011111110011011111011110000",
"10111011000000110011010010010100",
"01001100011111000110110110100110",
"00110010100000011100111110100101",
"01000100000110100111000100001000",
"00111010110101000010101111000001",
"11101000110100001011010101000000",
"10010110000111010000000100001001",
"11000100000111110010010111010101",
"10111010110011011110010110001101",
"01011010011011101101001110101010",
"00100100100010010011010000111011",
"11011110011010011001001010110100",
"10100000100011000100101001000111",
"11101001010101101110100100100110",
"10010101100110000111100011111101",
"00001011110100010011000000010011",
"01110011000111001010010011011001",
"10111001110111000001001010000110",
"11000101000101001110010110000000",
"01001011011010100001100110000101",
"00110011100010111111100101111101",
"11001111011000000010001001101101",
"10101111100100100011001010101101",
"10111100011011110011110110100110",
"11000010100010001111011101110011",
"00101010001100101010111010110010",
"01010100101101110110001100000111",
"01001001101001011101000101011000",
"00110101010001011001110101010011",
"10100100000110101001011100111101",
"11011010110100111111011101010001",
"10001001010110101111100101011011",
"11110101100101011010010010110000",
"10100101110000100011100110011101",
"11011001001010001011011000100101",
"10001001101010101010001010000001",
"11110101010000000000100100101111",
"01000100101100101000100010101111",
"00111010001101111000101000010011",
"10000010000010000001001111000010",
"11111100111100001100110111110101",
"00111101111100111110001010100110",
"01000001000001100101101110110100",
"00000001011011010010001111011100",
"01111101100010100010111000010000",
"10010111001100110110011110110010",
"11100111101101101010010111101100",
"00001001011000101111101001001000",
"01110101100100000101110111011011",
"11011100000011100100010000100100",
"10100010111001100101010000101110",
"00011000001111001110001111111100",
"01100110101011010111100111100010",
"00101000011010100000000001001110",
"01010110100011000000100010010010",
"00100001110010111011001011111001",
"01011101001000001101110101011110",
"10011010011001100110010010001011",
"11100100100011100011101000001001",
"01000010011000010001110001011100",
"00111100100100011001000001011011",
"11111001000100010001010010011010",
"10000101111000011101110001100001",
"00101111000110000000000010101011",
"01001111110101111001001101000011",
"00011001001100011000000000011011",
"01100101101110001001101110100111",
"00101101011001100011110100010101",
"01010001100011100101001001101001",
"00000110100011000110101110000010",
"01111000011010010101101101101110",
"01111101000001010110010100100011",
"00000001111101011010010101110010",
"00001111110111111111011101001110",
"01101111000100100100111011010011",
"01101011110010110001100111110100",
"00010011001000010101011010010001",
"00001011101100001101110011101111",
"01110011001110010100010111111001",
"01111000001000101101100100111000",
"00000110110010010011011110111010",
"11001001111110110010100000001001",
"10110101000000100111011111110000",
"10010011001011011000011110100110",
"11101011101111001101010100000000",
"11100101000010111101111011010111",
"10011001111010100100011000011110",
"01000101000000011101011101010111",
"00111001111111000101111010110000",
"10100000011010101011111011110000",
"11011110100010111001011011011010",
"10111101111100110011111100101010",
"11000001000001101011011000000001",
"11010011000111110000100101101010",
"10101011110011100000101001010111",
"10111000010011110010000111000011",
"11000110100111100011001011100000",
"00100101110011011110001100000001",
"01011001000111110010011111001101",
"11001010001101001001001001001111",
"10110100101101010111011111100000",
"10010101001000111010111110110000",
"11101001110010000011000000010101",
"11110000110110101001110010101011",
"10001110000101011110010000100010",
"11000101101011001000000001110011",
"10111001001111011111010100011110",
"01001100000101110000010111111111",
"00110010110110001111100100010100",
"01010001110100111100101011011011",
"00101101000110101011011110110001",
"00111001000111000111111001110110",
"01000101110100010110001101100011",
"01010100100110011001110001101101",
"00101010010101010101000101101001",
"00001110001101000001101100111011",
"01110000101101011110111111011011",
"00000001010000110100000010111011",
"01111101101001111101001011001011",
"00111001000101111011111010100111",
"01000101110101111111000100001100",
"11011010100110001110011001000101",
"10100100010101100100111110001011",
"00111011001010011101001100110111",
"01000011110000001111001110010110",
"01100100000101100011110110100111",
"00011010110110100001101001101001",
"00011010000010000111100100110101",
"01100100111100000001101011110100",
"11011001001011100101001111010010",
"10100101101110111111011111010111",
"10110110001111100110111100101100",
"11001000101011000001000111100011",
"10101011011101110000001011111000",
"11010011100001001010100001100010",
"10010011010101011010101010000010",
"11101011100110010101110001011111",
"10000011101111101100001001110111",
"11111011001010111100011011000001",
"01000010100000001110000011001101",
"00111100011111100100000101110110",
"00100011101001101000111110111001",
"01011011010001001011101101110100",
"01110001011000011000000000110111",
"00001101100100010100111111100110",
"01000111111001110110010101100000",
"00110111000011011001110000101101",
"00110001111001011010011101101011",
"01001101000011101010111100101001",
"01010010110010111000111000000101",
"00101100001000001111101010010010",
"01101010110110001010010111001000",
"00010100000101110100000000010000",
"11100010000010000110001111100011",
"10011100111100000100000001111100",
"01011011000111000110001111111010",
"00100011110100011000011011011001",
"00011001011110110110110111111001",
"01100101100000100101001110100110",
"11010000000000101100001000110011",
"10101110111110101001100101100110",
"11011001011000011110100010110101",
"10100101100100010000110010101111",
"11100000111110111100010101001110",
"10011110000000100010011001110001",
"00101101010110100011110100110110",
"01010001100101100010010110110010",
"11110101111111000110111100011000",
"10001001000000011100111011100111",
"11010011101111100010000001010010",
"10101011001011000101100101000000",
"10000110101010111000110100000000",
"11111000001111110000001010110000",
"10110100000110101010111100101001",
"11001010110100111101011010001001",
"01101111101001001101110000110010",
"00001111010001101100001100101110",
"11110111101000101010100010101001",
"10000111010010010111001111001100",
"01000101001011001011101010100110",
"00111001101111011011010100011101",
"00001100100001111110100110101111",
"01110010011100010001100010000001",
"01110111110100101010101011111001",
"00000111000110111000101100011110",
"11010110000001111101100101101101",
"10101000111100010011010101011011",
"00110100101011101110111100011101",
"01001010001110110101000011111010",
"01001000000100111110110000100011",
"00110110110111011000010110000100",
"01100010001011010000100100110001",
"00011100101111010101111100000001",
"00001010111100101110001010101111",
"01110100000001101110100101001100",
"10100110010011101100000010000101",
"11011000100111100111110101001000",
"10110111011110100011111001010000",
"11000111100000101111000111001011",
"01101001011001100001111110010011",
"00010101100011100110010010101001",
"11010100110010000111111110000011",
"10101010001000110110111011011000",
"00000010100111010000111010101110",
"01111100010100001010001100011110",
"01101000000111101011100111001010",
"00010110110011100111000110110100",
"10000100111001010100001100110110",
"11111010000011101110110110000111",
"00010011110011000110111001111101",
"01101011001000000100100111010000",
"00101010001011111001100100100010",
"01010100101110101001101110011101",
"11111010000101110101111001001010",
"10000100110110000111101010000101",
"10001110111001001010010110111110",
"11110000000011110100111111110110",
"11110100111100010101001100001110",
"10001010000001111100100010110101",
"00111111101000100111111100011101",
"00111111010010011010011101001110",
"11001000010001010100011000101011",
"10110110101001100001101010011010",
"01011110011110110001010000001010",
"00100000100000101000001001010100",
"01100100111110000101011011001111",
"00011010000000111111001011011000",
"10001011100001010100100011000000",
"11110011011101011101100111000011",
"10100001000101010000010000101101",
"11011101110110111110010100111000",
"00100111101010101111001111000010",
"01010111001111111010110111101001",
"01100100111111010001010011100110",
"00011010000000010111100111011100",
"10011100100010011110110101010000",
"11100010011011011001001100110000",
"10101100110111010011000100100011",
"11010010000101000010010010010001",
"11001101101101111111001101110000",
"10110001001100100010001001101100",
"01010000101010101011001111111001",
"00101110001111111111010110001000",
"11111001000011110000111001100000",
"10000101111001010000111010010010",
"10010111111011101000100101110010",
"11100111000010010101111011101100",
"10100011001000101110111010010011",
"11011011110010010001110101011010",
"00101011000001011010000010100001",
"01010011111101010011100000010101",
"11111001011000001001000011011110",
"10000101100100011110101011000110",
"10111110101000000101110110011001",
"11000000010011000101010101000101",
"10001110010010101000100100111011",
"11110000101000011100100111011010",
"11111010110010110111110011001101",
"10000100001000010000100000110001",
"10111111000100010000111010101100",
"10111111111000011110010110011101",
"00100101001111010001000100011001",
"01011001101011010101000001111110",
"01001100101111100111001011111111",
"00110010001011000000111001101111",
"11110001001010011111001001000010",
"10001101110000001101000001010111",
"10100111101000111011100100001010",
"11010111010010000010010010100110",
"00011001100111101011110000011100",
"01100101010011100110111010101111",
"11110101000100111110110110101011",
"10001001110111011000001100111001",
"10111101001010101111111000110100",
"11000001101111111010001000110011",
"01001001110110001100100111001100",
"00110101000101110010011011101111",
"11011100001000110101110101111010",
"10100010110010001001010011010011",
"10101100101010101001000000110110",
"11010010010000000001110111001000",
"01011000011000111110110100011110",
"00100110100011111100010000001100",
"10010000101010011011001011000111",
"11101110010000010001100001110111",
"00000100011001000000100011000010",
"01111010100011111011001010011111",
"11100001001010011111000100010000",
"10011101110000001101000110110010",
"01001110010100111100100101101011",
"00110000100110101011100010111110",
"10100001101001011111011000011110",
"11011101010001010111000110001010",
"11000100010010010010001101001110",
"10111010101000101110100111000001",
"00010111100011101001110111111011",
"01100111011001011100001100010110",
"11010111101011001100100101101100",
"10100111001111011010010011100101",
"01010011011110100011100011110101",
"00101011100000101111010010011001",
"00110100100011100000001101111111",
"01001010011001101011110100000110",
"01011011100101001111010110011101",
"00100011010110111111101010111000",
"10110110101100010010001010101100",
"11001000001110001111110100000111",
"01000110110100101000100101011010",
"00111000000110111010001111110100",
"00010010011010010111011111001001",
"01101100100011000101101001110100",
"10011001111111010111111001000010",
"11100101000000010100010000001011",
"10011001100010000011101010100101",
"11100101011100001000100100111000",
"10000001110100011010111110011110",
"11111101000111000100010110010010",
"01001001100110110110110100001011",
"00110101010100101101001110111100",
"10011101000110111100100011110110",
"11100001110100100101011101010111",
"00000011001101101010000001101010",
"01111011101100110110110100011011",
"00001011100000000001000011111100",
"01110011011111111101111000001101",
"10101101001001100010100000110001",
"11010001110001010011011000001001",
"11111100111100101101100101001000",
"10000010000001101110111010000101",
"11100010010000010000010111111101",
"10011100101010011100001100000110",
"01110110000111100111011100100101",
"00001000110011101100100010000110",
"00011000111110110011100011011110",
"01100110000000100110111100110011",
"00001000100010000000101100110000",
"01110110011100001101110100100001",
"11110111001000010010110000101011",
"10000111110010110100111101100001",
"01100010100000001101101110110000",
"00011100011111100100101110001101",
"01000010110101111010111000011011",
"00111100000101111110110111000000",
"01110100010110000000100011011011",
"00001010100101111010110111101110",
"10100111001001011000101011111011",
"11010111110001011111000101010010",
"11111010010011000010110000100111",
"10000100101000000111110111100100",
"11011001001001010101100100100111",
"10100101110001100010110011111001",
"10001000101100000010111001111110",
"11110110001110011111110101101010",
"01010110001010011011010000110001",
"00101000110000010001011011011100",
"00100011110110111011110101001001",
"01011011000101010001111101000010",
"10110111001111101110111001110001",
"11000111101010111001111100110001",
"00001000001000101100110111111111",
"01110110110010010100010110011001",
"01110001001110111010100011001111",
"00001101101011101001110100111101",
"10110000010011101111110111101011",
"11001110100111100100111001000101",
"11001111111101001011000111100110",
"10101111000001011110100111101000",
"01011001111000110011110100110111",
"00100101000100000011001101010101",
"10001000001100011001110110100110",
"11110110101110000111110011110011",
"01010000101000001000001000000110",
"00101110010011000010011011100110",
"00111000111000100111001011011010",
"01000110000100001011010000110010",
"10100111011010010011010010000010",
"11010111100011001000001011110010",
"00111011001000100100001101011011",
"01000011110010011111000110010001",
"11010000110010001111010111011100",
"10101110001000110000111010011000",
"00111001000111010101010111000111",
"01000101110100000100010011010110",
"11110000101000111001011000010100",
"10001110010010000100111101101100",
"01101101101010010110001111010100",
"00010001010000010111001001110111",
"00010010100101101110011001011011",
"01101100010110010010011010010011",
"10110101010011011110100111101111",
"11001001100111110010001001110010",
"00111110011010000100011010110100",
"01000000100011010001001011001101",
"10011000111110101111100101111111",
"11100110000000101001000000100010",
"00110000110000000111010001101011",
"01001110001010100100001101101110",
"00100111100011100100110110111011",
"01010111011001100100010010101000",
"10110000000001011000100101111000",
"11001110111101010110001010011100",
"01000111000001111100101010001010",
"00110111111100010100111111001101",
"01111010110010010011011100100011",
"00000100001000101101100110110010",
"01000101100111101001011001100000",
"00111001010011101001111111001110",
"01011111111100100011101100111001",
"00011111000001110100011010010001",
"01000011111001111100110001010000",
"00111011000011010101110101001010",
"10010101000010000111011000111111",
"11101001111100000010000000101010",
"10001010001101000101010101110000",
"11110100101101011011010100100001",
"10001100010011000010110000010000",
"11110010101000000111110111110110",
"00011010001010110101111110110001",
"01100100101111110011010100110000",
"10011100110001100000101110001011",
"11100010001001010111010100010000",
"10111001100111001100011011000111",
"11000101010100010000001011001110",
"01110110000000101101110001011111",
"00001000111110100110011101001000",
"11001001111001011001011011011111",
"10110101000011101011100101110010",
"00111011100001110110101110101100",
"01000011011100011111100011011001",
"00110001011001110000001001101101",
"01001101100011011101100011010101",
"10100001001100111100111111111011",
"11011101101101100011101111111110",
"11101100001100110000000010100011",
"10010010101101110000111100010101",
"11111000010110010000101001011011",
"10000110100101101111100111111010",
"10111110001011110111001011000101",
"11000000101110101100010001101011",
"10110010100100100111000010111111",
"11001100010111111100001101101100",
"00001001000001100111011010101011",
"01110101111100111011000110111110",
"11001101010001101111001101010010",
"10110001101001001011010001001110",
"10001011000110001000010101100000",
"11110011110101101101011110110001",
"10101010010010111001111110101001",
"11010100101000001110110010100000",
"00110110111010111001110010100100",
"01001000000010110001001110000001",
"00000011000011001110001100101011",
"01111011111010001001010100111100",
"00110110100000000010011010110110",
"01001000011111111011001010101011",
"11010011101100011100100111001111",
"10101011001110000100111100100000",
"00111110011001100101111010100100",
"01000000100011100011110110101110",
"11011101100101001000011110000111",
"10100001010111001001110111000011",
"01111101100001111001100100110100",
"00000001011100011010011110011001",
"11111011100101110011010110111110",
"10000011010110001011010010010001",
"11111011100110010001111100101110",
"10000011010101011111111111100100",
"11001110001010111110100100100100",
"10110000101111101001110001001111",
"10111011110111011110011110011000",
"11000011000100111010101011000010",
"11110101110001100111011011101100",
"10001001001001010001101110001010",
"01101010011011010010101111101011",
"00010100100010100010100101011110",
"11000110011000101101011000000010",
"10111000100100000111010011110001",
"10101010011111111011110101000001",
"11010100100000000010000101101000",
"00011101011001000100001000110111",
"01100001100011111000111001110011",
"01010100100101101101110000011011",
"00101010010110010011010101010100",
"10001110010110011101001011101010",
"11110000100101100110111011110111");

  signal op,ans1,ans,answ,low,high: std_logic_vector(31 downto 0);
  signal addr: std_logic_vector(19 downto 0) := (others=>'0');
  signal miss: std_logic_vector(31 downto 0) := (others=>'0');
  signal rom_o: std_logic_vector(7 downto 0) := (others=>'1');
  signal uart_go: std_logic;
  signal uart_busy: std_logic := '0';
  signal iter: std_logic_vector(31 downto 0) := (others=>'0');
  signal state: std_logic_vector(4 downto 0) := (others=>'0');
  signal state2: std_logic_vector(4 downto 0) := (others=>'0');

begin

  ib: IBUFG port map (
   i=>MCLK1,
   o=>iclk);
  bg: BUFG port map (
    i=>iclk,
    o=>clk);

  finver:finv port map
    (clk, op, ans);

  rs232c: u232c generic map (wtime=>x"1ADB")
  port map (
    clk=>clk,
    data=>rom_o,
    go=>uart_go,
    busy=>uart_busy,
    tx=>rs_tx);


 cal: process(clk)
 begin
   if rising_edge(clk) then-- hoge clk後に返答
     if state = "00000" and addr = 3944 then -- 最後はnop
       state<="00000";
     elsif state = "00000" then
       state<=state+1;
       addr<=addr+2;
       op<=rom(conv_integer(addr));
       ans1<=rom(conv_integer(addr+1));
     elsif state = "00001" then
       state<=state+1;
     elsif state = "00010" then
       state<=state+1;
       answ<=ans;
       state2<="00000";
     elsif state = "00011" and uart_go = '1'then --op1の出力
       state2<=state2+1;
       if op(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "00100" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "00101" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "00110" and uart_go = '1'then --op2の出力
       --state2<=state2+1;
       --if op2(31-conv_integer(state2)) = '1' then
         --rom_o<=x"31";
       --else
         --rom_o<=x"30";
       --end if;
       --if state2 = "11111" then
         state<=state+1;
         --state2<="00000";
       --end if;
     elsif state = "00111" and uart_go = '1'then -- 改行
       state<=state+1;
       --rom_o<=x"0d";
     elsif state = "01000" and uart_go = '1'then
       state<=state+1;
       --rom_o<=x"0a";
     elsif state = "01001" and uart_go = '1'then --outputの出力
       state2<=state2+1;
       if answ(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01010" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01011" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01100" and uart_go = '1'then --answerの出力
       state2<=state2+1;
       if ans1(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01101" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01110" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01111" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10000" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10001" then --low,highとの比較
       state<=state+1;
       low<=ans1 - 5;
     elsif state = "10010" then
       state<=state+1;
       high<=ans1 + 5;
     elsif state = "10011" then
       iter<=iter+1;
       state<=state+1;
       if high < answ or low > answ then
         miss<=miss+1;
       end if;
     elsif state = "10100" and uart_go = '1'then --iterの出力
       state2<=state2+1;
       if iter(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "10101" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10110" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10111" and uart_go = '1'then --missの出力
       state2<=state2+1;
       if miss(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "11000" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11001" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "11010" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11011" and uart_go = '1'then
       state<="00000";
       rom_o<=x"0a";
     end if;
   end if;
 end process;

    send_msg: process(clk)
  begin
    if rising_edge(clk) then
      if uart_busy='0' and uart_go='0' then
        uart_go<='1';
      else
        uart_go<='0';
      end if;
    end if;
  end process;
  
end VHDL;
