library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity blockram2 is

  generic (
    dwidth : integer := 13;
    awidth : integer := 10);

  port (
    clk  : in  std_logic;
    we   : in  std_logic;
    di   : in  std_logic_vector(dwidth - 1 downto 0);
    do   : out std_logic_vector(dwidth - 1 downto 0);
    addr : in  std_logic_vector(awidth - 1 downto 0));

end blockram2;

architecture behavioral of blockram2 is

  type ram_type is
    array(0 to (2 ** awidth) - 1) of std_logic_vector(dwidth - 1 downto 0);

  signal ram : ram_type := (
"0110100111100",
"0110100110000",
"0110100100100",
"0110100011010",
"0110100001111",
"0110100000011",
"0110011111000",
"0110011101110",
"0110011100001",
"0110011011000",
"0110011001100",
"0110011000000",
"0110010110101",
"0110010101100",
"0110010100000",
"0110010010110",
"0110010001011",
"0110010000000",
"0110001110101",
"0110001101011",
"0110001100000",
"0110001010101",
"0110001001011",
"0110001000000",
"0110000110100",
"0110000100110",
"0110000011110",
"0110000010011",
"0110000001100",
"0110000000000",
"0101111110101",
"0101111101100",
"0101111100010",
"0101111011000",
"0101111001101",
"0101111000010",
"0101110111000",
"0101110110000",
"0101110100100",
"0101110011011",
"0101110010000",
"0101110000111",
"0101101111100",
"0101101101111",
"0101101100111",
"0101101011110",
"0101101010100",
"0101101001001",
"0101101000000",
"0101100110110",
"0101100101101",
"0101100100011",
"0101100011001",
"0101100001101",
"0101100000110",
"0101011111011",
"0101011110011",
"0101011101001",
"0101011100000",
"0101011010101",
"0101011001100",
"0101011000011",
"0101010111000",
"0101010101110",
"0101010100100",
"0101010011010",
"0101010010011",
"0101010001010",
"0101010000000",
"0101001110110",
"0101001101101",
"0101001100100",
"0101001011011",
"0101001010000",
"0101001001000",
"0101000111110",
"0101000110101",
"0101000101100",
"0101000100100",
"0101000011010",
"0101000010010",
"0101000001000",
"0100111111110",
"0100111110101",
"0100111101101",
"0100111100100",
"0100111011010",
"0100111010010",
"0100111001001",
"0100111000000",
"0100110111000",
"0100110101110",
"0100110100111",
"0100110011100",
"0100110010100",
"0100110001100",
"0100110000011",
"0100101111010",
"0100101110001",
"0100101101001",
"0100101100000",
"0100101011000",
"0100101010000",
"0100101000110",
"0100100111110",
"0100100110101",
"0100100101100",
"0100100100011",
"0100100011011",
"0100100010100",
"0100100001010",
"0100100000011",
"0100011111001",
"0100011110010",
"0100011101001",
"0100011100000",
"0100011011000",
"0100011001111",
"0100011000111",
"0100010111110",
"0100010110111",
"0100010101100",
"0100010100110",
"0100010011111",
"0100010010110",
"0100010001110",
"0100010000110",
"0100001111110",
"0100001110110",
"0100001101110",
"0100001100110",
"0100001011110",
"0100001010100",
"0100001001101",
"0100001000101",
"0100000111111",
"0100000110101",
"0100000101111",
"0100000100101",
"0100000011110",
"0100000010110",
"0100000001111",
"0100000000110",
"0100000000000",
"0011111110111",
"0011111101110",
"0011111101000",
"0011111100000",
"0011111011000",
"0011111010000",
"0011111001001",
"0011111000000",
"0011110111001",
"0011110110001",
"0011110101001",
"0011110100010",
"0011110011001",
"0011110010011",
"0011110001100",
"0011110000100",
"0011101111100",
"0011101110100",
"0011101101110",
"0011101100110",
"0011101011111",
"0011101010111",
"0011101010000",
"0011101001000",
"0011101000000",
"0011100111010",
"0011100110010",
"0011100101011",
"0011100100100",
"0011100011100",
"0011100010101",
"0011100001110",
"0011100000110",
"0011011111110",
"0011011110111",
"0011011110000",
"0011011101010",
"0011011100010",
"0011011011011",
"0011011010011",
"0011011001100",
"0011011000110",
"0011010111111",
"0011010110111",
"0011010110001",
"0011010101001",
"0011010100010",
"0011010011011",
"0011010010001",
"0011010001110",
"0011010000110",
"0011010000000",
"0011001111000",
"0011001110001",
"0011001101010",
"0011001100100",
"0011001011100",
"0011001010111",
"0011001001110",
"0011001001001",
"0011001000000",
"0011000111010",
"0011000110100",
"0011000101101",
"0011000100110",
"0011000011111",
"0011000011000",
"0011000010010",
"0011000001011",
"0011000000100",
"0010111111100",
"0010111110111",
"0010111110000",
"0010111101010",
"0010111100011",
"0010111011100",
"0010111010110",
"0010111001111",
"0010111001001",
"0010111000001",
"0010110111011",
"0010110110101",
"0010110101110",
"0010110101000",
"0010110100000",
"0010110011010",
"0010110010011",
"0010110001101",
"0010110001000",
"0010110000000",
"0010101111010",
"0010101110100",
"0010101101110",
"0010101100111",
"0010101100001",
"0010101011011",
"0010101010100",
"0010101001110",
"0010101000111",
"0010101000000",
"0010100111100",
"0010100110011",
"0010100101110",
"0010100101000",
"0010100100010",
"0010100011100",
"0010100010110",
"0010100001111",
"0010100001001",
"0010100000010",
"0010011111101",
"0010011110110",
"0010011101111",
"0010011101011",
"0010011100101",
"0010011011101",
"0010011010110",
"0010011010001",
"0010011001001",
"0010011000101",
"0010011000000",
"0010010111001",
"0010010110011",
"0010010101110",
"0010010100110",
"0010010100000",
"0010010011011",
"0010010010101",
"0010010001110",
"0010010001001",
"0010010000011",
"0010001111100",
"0010001110111",
"0010001110000",
"0010001101011",
"0010001100110",
"0010001100000",
"0010001011010",
"0010001010100",
"0010001001111",
"0010001001000",
"0010001000011",
"0010000111100",
"0010000110110",
"0010000110000",
"0010000101011",
"0010000100110",
"0010000100000",
"0010000011010",
"0010000010011",
"0010000001110",
"0010000001000",
"0010000000100",
"0001111111101",
"0001111111000",
"0001111110010",
"0001111101101",
"0001111100111",
"0001111100001",
"0001111011100",
"0001111010101",
"0001111010000",
"0001111001011",
"0001111000101",
"0001110111110",
"0001110111010",
"0001110110100",
"0001110101110",
"0001110101000",
"0001110100011",
"0001110011110",
"0001110011001",
"0001110010011",
"0001110001110",
"0001110001000",
"0001110000100",
"0001101111100",
"0001101111001",
"0001101110010",
"0001101101101",
"0001101101000",
"0001101100010",
"0001101011101",
"0001101011000",
"0001101010010",
"0001101001100",
"0001101000111",
"0001101000010",
"0001100111100",
"0001100110111",
"0001100110010",
"0001100101100",
"0001100100111",
"0001100100010",
"0001100011101",
"0001100010111",
"0001100010001",
"0001100001100",
"0001100000110",
"0001100000011",
"0001011111110",
"0001011111000",
"0001011110010",
"0001011101101",
"0001011101001",
"0001011100100",
"0001011011110",
"0001011011001",
"0001011010011",
"0001011001100",
"0001011001001",
"0001011000101",
"0001010111111",
"0001010111000",
"0001010110101",
"0001010101111",
"0001010101010",
"0001010100110",
"0001010100000",
"0001010011011",
"0001010010101",
"0001010010010",
"0001010001100",
"0001010001000",
"0001010000000",
"0001001111101",
"0001001110111",
"0001001110100",
"0001001101110",
"0001001101010",
"0001001100010",
"0001001011111",
"0001001011011",
"0001001010101",
"0001001010001",
"0001001001011",
"0001001000110",
"0001001000010",
"0001000111101",
"0001000111000",
"0001000110011",
"0001000101110",
"0001000101000",
"0001000100100",
"0001000100000",
"0001000011011",
"0001000010110",
"0001000010001",
"0001000001100",
"0001000000101",
"0001000000010",
"0001000000000",
"0000111111000",
"0000111110101",
"0000111101111",
"0000111101010",
"0000111100101",
"0000111100010",
"0000111011100",
"0000111011000",
"0000111010011",
"0000111001110",
"0000111001010",
"0000111000101",
"0000111000000",
"0000110111100",
"0000110110111",
"0000110110010",
"0000110101101",
"0000110101000",
"0000110100011",
"0000110100000",
"0000110011011",
"0000110010110",
"0000110010010",
"0000110001101",
"0000110001001",
"0000110000101",
"0000110000000",
"0000101111010",
"0000101110101",
"0000101110001",
"0000101101101",
"0000101101001",
"0000101100101",
"0000101100000",
"0000101011010",
"0000101010101",
"0000101010010",
"0000101001101",
"0000101001001",
"0000101000100",
"0000101000000",
"0000100111011",
"0000100110111",
"0000100110010",
"0000100101110",
"0000100101001",
"0000100100100",
"0000100100001",
"0000100011100",
"0000100011000",
"0000100010100",
"0000100001111",
"0000100001010",
"0000100000110",
"0000100000000",
"0000011111100",
"0000011111001",
"0000011110100",
"0000011101111",
"0000011101011",
"0000011101000",
"0000011100011",
"0000011011110",
"0000011011011",
"0000011010110",
"0000011010010",
"0000011001101",
"0000011001001",
"0000011000101",
"0000011000000",
"0000010111100",
"0000010111000",
"0000010110011",
"0000010101111",
"0000010101011",
"0000010100111",
"0000010100011",
"0000010011110",
"0000010011001",
"0000010010101",
"0000010010001",
"0000010001100",
"0000010001001",
"0000010000110",
"0000010000000",
"0000001111101",
"0000001111000",
"0000001110011",
"0000001110000",
"0000001101100",
"0000001101000",
"0000001100011",
"0000001100000",
"0000001011010",
"0000001010111",
"0000001010011",
"0000001001110",
"0000001001010",
"0000001000111",
"0000001000011",
"0000000111101",
"0000000111010",
"0000000110111",
"0000000110010",
"0000000101111",
"0000000101011",
"0000000100110",
"0000000100010",
"0000000011111",
"0000000011011",
"0000000010101",
"0000000010001",
"0000000001101",
"0000000001001",
"0000000000101",
"0000000000000",
"1111111111111",
"1111111101000",
"1111111011000",
"1111111001000",
"1111110111001",
"1111110101010",
"1111110011000",
"1111110001010",
"1111101111010",
"1111101101010",
"1111101011010",
"1111101001011",
"1111100111010",
"1111100101110",
"1111100011110",
"1111100001101",
"1111100000000",
"1111011101110",
"1111011100001",
"1111011010001",
"1111011000011",
"1111010110011",
"1111010100101",
"1111010010101",
"1111010000111",
"1111001111010",
"1111001101000",
"1111001011001",
"1111001001010",
"1111000111011",
"1111000101101",
"1111000011110",
"1111000001111",
"1111000000000",
"1110111110001",
"1110111100101",
"1110111010110",
"1110111001000",
"1110110111000",
"1110110101011",
"1110110011101",
"1110110001111",
"1110110000000",
"1110101110001",
"1110101100011",
"1110101010100",
"1110101000111",
"1110100111010",
"1110100101101",
"1110100011100",
"1110100010000",
"1110100000000",
"1110011110011",
"1110011100110",
"1110011011001",
"1110011001011",
"1110010111110",
"1110010110001",
"1110010100001",
"1110010010010",
"1110010000111",
"1110001111000",
"1110001101011",
"1110001011110",
"1110001010000",
"1110001000010",
"1110000110101",
"1110000100111",
"1110000011010",
"1110000001110",
"1110000000000",
"1101111110010",
"1101111100111",
"1101111011001",
"1101111001100",
"1101110111111",
"1101110110011",
"1101110100110",
"1101110011000",
"1101110001011",
"1101101111110",
"1101101110010",
"1101101100110",
"1101101011000",
"1101101001011",
"1101101000000",
"1101100110001",
"1101100100100",
"1101100011001",
"1101100001010",
"1101011111111",
"1101011110001",
"1101011100110",
"1101011011011",
"1101011001110",
"1101011000000",
"1101010110011",
"1101010101000",
"1101010011100",
"1101010010000",
"1101010000011",
"1101001111000",
"1101001101011",
"1101001100000",
"1101001010011",
"1101001001000",
"1101000111010",
"1101000101111",
"1101000100001",
"1101000010110",
"1101000001100",
"1100111111111",
"1100111110001",
"1100111100111",
"1100111011101",
"1100111010000",
"1100111000011",
"1100110110111",
"1100110101011",
"1100110100001",
"1100110010101",
"1100110001011",
"1100101111111",
"1100101110011",
"1100101100111",
"1100101011001",
"1100101001111",
"1100101000101",
"1100100110111",
"1100100101101",
"1100100100011",
"1100100010111",
"1100100001011",
"1100100000000",
"1100011110101",
"1100011101010",
"1100011011111",
"1100011010010",
"1100011001000",
"1100010111100",
"1100010110001",
"1100010100101",
"1100010011010",
"1100010010000",
"1100010000101",
"1100001111010",
"1100001101110",
"1100001100101",
"1100001011010",
"1100001001101",
"1100001000011",
"1100000111010",
"1100000101100",
"1100000100001",
"1100000010111",
"1100000001100",
"1100000000010",
"1011111111000",
"1011111101101",
"1011111100100",
"1011111010110",
"1011111001111",
"1011111000011",
"1011110111001",
"1011110101110",
"1011110100011",
"1011110010111",
"1011110001101",
"1011110000100",
"1011101111000",
"1011101110000",
"1011101100110",
"1011101011001",
"1011101001110",
"1011101000111",
"1011100111011",
"1011100101111",
"1011100100111",
"1011100011100",
"1011100010010",
"1011100001000",
"1011011111111",
"1011011110100",
"1011011101001",
"1011011011110",
"1011011010110",
"1011011001011",
"1011011000011",
"1011010110111",
"1011010101100",
"1011010100100",
"1011010011000",
"1011010010001",
"1011010000101",
"1011001111100",
"1011001110001",
"1011001100111",
"1011001011101",
"1011001010011",
"1011001001001",
"1011001000000",
"1011000111000",
"1011000101110",
"1011000100100",
"1011000011010",
"1011000010000",
"1011000000111",
"1010111111100",
"1010111110100",
"1010111101001",
"1010111011111",
"1010111010110",
"1010111001110",
"1010111000011",
"1010110111001",
"1010110110000",
"1010110101000",
"1010110011101",
"1010110010011",
"1010110001011",
"1010110000000",
"1010101111000",
"1010101101111",
"1010101101000",
"1010101011110",
"1010101010010",
"1010101001011",
"1010101000010",
"1010100111000",
"1010100101100",
"1010100100100",
"1010100011101",
"1010100010100",
"1010100001001",
"1010100000000",
"1010011111001",
"1010011101111",
"1010011100111",
"1010011011101",
"1010011010101",
"1010011001011",
"1010011000011",
"1010010111001",
"1010010110000",
"1010010101000",
"1010010011110",
"1010010010011",
"1010010001100",
"1010010000011",
"1010001111011",
"1010001110011",
"1010001101001",
"1010001100010",
"1010001011001",
"1010001001111",
"1010001000111",
"1010000111110",
"1010000110011",
"1010000101011",
"1010000100010",
"1010000011010",
"1010000010000",
"1010000001001",
"1010000000000",
"1001111110111",
"1001111101110",
"1001111101001",
"1001111011110",
"1001111010110",
"1001111001101",
"1001111000100",
"1001110111101",
"1001110110010",
"1001110101010",
"1001110100011",
"1001110011010",
"1001110010011",
"1001110001010",
"1001110000000",
"1001101111000",
"1001101110010",
"1001101101000",
"1001101100000",
"1001101011001",
"1001101010001",
"1001101001001",
"1001101000000",
"1001100110111",
"1001100101101",
"1001100100111",
"1001100011101",
"1001100010110",
"1001100001111",
"1001100000111",
"1001011111110",
"1001011110110",
"1001011101110",
"1001011101000",
"1001011011110",
"1001011010110",
"1001011001110",
"1001011000110",
"1001010111110",
"1001010110110",
"1001010101110",
"1001010100110",
"1001010011110",
"1001010010111",
"1001010001110",
"1001010000101",
"1001001111111",
"1001001110101",
"1001001101110",
"1001001101000",
"1001001011111",
"1001001010110",
"1001001010001",
"1001001001000",
"1001001000000",
"1001000111001",
"1001000101111",
"1001000101000",
"1001000011111",
"1001000011010",
"1001000010001",
"1001000001010",
"1001000000011",
"1000111111010",
"1000111110101",
"1000111101100",
"1000111100100",
"1000111011101",
"1000111010100",
"1000111001110",
"1000111000101",
"1000110111110",
"1000110110111",
"1000110101110",
"1000110100110",
"1000110011111",
"1000110011000",
"1000110010000",
"1000110001010",
"1000110000100",
"1000101111100",
"1000101110100",
"1000101101100",
"1000101100110",
"1000101011110",
"1000101010110",
"1000101010000",
"1000101001000",
"1000101000000",
"1000100111001",
"1000100110010",
"1000100101011",
"1000100100010",
"1000100011100",
"1000100010100",
"1000100001110",
"1000100000111",
"1000100000000",
"1000011111000",
"1000011110001",
"1000011101001",
"1000011100010",
"1000011011100",
"1000011010101",
"1000011010000",
"1000011000111",
"1000011000000",
"1000010111001",
"1000010110000",
"1000010101011",
"1000010100011",
"1000010011100",
"1000010010101",
"1000010001101",
"1000010000111",
"1000010000000",
"1000001111001",
"1000001110001",
"1000001101011",
"1000001100011",
"1000001011101",
"1000001010101",
"1000001010000",
"1000001001001",
"1000001000000",
"1000000111010",
"1000000110101",
"1000000101100",
"1000000100111",
"1000000100000",
"1000000010111",
"1000000010010",
"1000000001100",
"1000000000101",
"0111111111110",
"0111111110111",
"0111111101111",
"0111111101010",
"0111111100011",
"0111111011011",
"0111111010101",
"0111111001110",
"0111111001001",
"0111111000000",
"0111110111001",
"0111110110100",
"0111110101110",
"0111110101000",
"0111110100000",
"0111110011010",
"0111110010001",
"0111110001101",
"0111110000101",
"0111110000000",
"0111101111001",
"0111101110010",
"0111101101100",
"0111101100110",
"0111101011111",
"0111101011000",
"0111101010011",
"0111101001101",
"0111101000110",
"0111100111111",
"0111100110111",
"0111100110001",
"0111100101011",
"0111100100100",
"0111100011101",
"0111100011000",
"0111100010010",
"0111100001100",
"0111100000101",
"0111100000000",
"0111011111000",
"0111011110011",
"0111011101101",
"0111011100111",
"0111011100000",
"0111011011001",
"0111011010010",
"0111011001101",
"0111011000101",
"0111011000000",
"0111010111010",
"0111010110011",
"0111010101101",
"0111010101010",
"0111010011111",
"0111010011011",
"0111010010011",
"0111010001110",
"0111010001001",
"0111010000000",
"0111001111101",
"0111001110111",
"0111001110001",
"0111001101011",
"0111001100101",
"0111001011110",
"0111001010111",
"0111001010001",
"0111001001010",
"0111001000100",
"0111000111111",
"0111000111000",
"0111000110010",
"0111000101101",
"0111000100110",
"0111000100000",
"0111000011011",
"0111000010100",
"0111000001110",
"0111000001001",
"0111000000011",
"0110111111101",
"0110111110111",
"0110111110000",
"0110111101010",
"0110111100111",
"0110111100000",
"0110111011011",
"0110111010101",
"0110111001100",
"0110111000111",
"0110111000010",
"0110110111101",
"0110110110101",
"0110110110000",
"0110110101010",
"0110110100110",
"0110110011111",
"0110110011001",
"0110110010011",
"0110110001101",
"0110110001000",
"0110110000011",
"0110101111101",
"0110101110110",
"0110101110010",
"0110101101011",
"0110101100110",
"0110101100000",
"0110101011011",
"0110101010100",
"0110101001111",
"0110101001001",
"0110101000011");

  signal reg_addr : std_logic_vector(awidth - 1 downto 0);

begin

  process(clk)
  begin
    if rising_edge(clk) then
      if we = '1' then
        ram(conv_integer(addr)) <= di;
      end if;
      reg_addr <= addr;
    end if;
  end process;

  do <= ram(conv_integer(reg_addr));

end behavioral;
