library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity fputop is
  port(MCLK1: in std_logic;
       RS_TX: out std_logic);
  end fputop;

architecture VHDL of fputop is

component fsqrt
  port(clk: in std_logic;
       op:  in std_logic_vector(31 downto 0);
       ans:       out std_logic_vector(31 downto 0) := x"00000000"
       );
end component;

component u232c
  generic (wtime: std_logic_vector(15 downto 0) := x"1ADB");
  Port ( clk  : in  STD_LOGIC;
         data : in  STD_LOGIC_VECTOR (7 downto 0);
         go   : in  STD_LOGIC;
         busy : out STD_LOGIC;
         tx   : out STD_LOGIC);
end component;

  signal clk,iclk: std_logic;
  type rom_t is array(0 to 3967) of std_logic_vector(31 downto 0);
  constant rom: rom_t := ("01001000111001000000111100100001",
"01000100001010101101101011111010",
"01101100110001100111001010111001",
"01010110000111110110000011000110",
"00110111000000010101000100101000",
"00111011001101011111001010111111",
"00001011100100010101011111001101",
"00100101100010000110010101100111",
"00100110101111110100010010111101",
"00110011000111000111011111101001",
"00010111111101111111010110110011",
"00101011101100100010011101101100",
"00010001111111111000000111110111",
"00101000101101001101100001011101",
"01100101011000101111011100111011",
"01010010011100010000101111001101",
"00001000000011001100011110001110",
"00100011101111011101011101000010",
"01101010101110111001011010001000",
"01010101000110101111010010100111",
"01010010011100000001000101100000",
"01001000111101111110011111101101",
"00010010101001011010111011110011",
"00101001000100011010000010111011",
"01110110101110111101011010100111",
"01011011000110110000111100100000",
"00110100010101100010101001000101",
"00111001111010100010011001101100",
"00100111001010110010110001000011",
"00110011010100010101010100111000",
"01010001101111111111010100011101",
"01001000100111001011111111111101",
"00001100111011010101110111101001",
"00100110001011100100111010011011",
"00101110101111000110101011000101",
"00110111000110110100110000110111",
"01001001101100100101111101100110",
"01000100100101110001101000000011",
"01010111011001101111010100101010",
"01001011011100110010100000011011",
"01101110001100000101010100001000",
"01010110110101000111011011010101",
"00110111011111001011110010010110",
"00111011011111100101110011110011",
"01011100001000011001001110111100",
"01001101110010110110000101111001",
"01000110011010000010111011111101",
"01000010111100111100110100010101",
"00111010111110010000100000011111",
"00111101001100101000100111100110",
"01111101111010010101111011101011",
"01011110101011001101010101100111",
"00100010001111100111111010000101",
"00110000110111001101010011011000",
"00010110101111100011000011111001",
"00101011000111000000011011110110",
"01001000100111010101111011011001",
"01000100000011011110110101110010",
"00000111101100101000100100010100",
"00100011100101110010101110101001",
"01011111101000100100000000011010",
"01001111100100000001110001111010",
"00110101011000111101000110010010",
"00111010011100010111111110100010",
"00111110101100111101101000111100",
"00111111000101111011101000100100",
"01101011001100111001011111100111",
"01010101010101100110101101111111",
"01011100001000110001011001001111",
"01001101110011000101010000110100",
"01010110101010111100111111101111",
"01001011000101000100110000000000",
"01111101001100110001100111011110",
"01011110010101100010000000110110",
"01000001100001100000110110001010",
"01000000100000101111110111010001",
"01011110101110001001011101111110",
"01001111000110011011011010010011",
"01100111111011101011000001100110",
"01010011101011101100101010110111",
"00010011111101100001111011101010",
"00101001101100010111110111111100",
"01110001010111100100011001110001",
"01011000011011101000101011010101",
"01011110101010101000011100001101",
"01001111000100111011110111001100",
"01001000010011000100100100101111",
"01000011111001001010111110001110",
"00011000100010010111001010110100",
"00101100000001001010001111010010",
"01011110101001101110011010110101",
"01001111000100100010100101111101",
"00011010000011000011111001001100",
"00101100101111010111101010100001",
"00100101011101101101000010011110",
"00110010011110110101110110010001",
"00001101011000110101000101111011",
"00100110011100010011101110110101",
"01100011101111101001110110110011",
"01010001100111000011001110001000",
"01111100110111011100010111001000",
"01011110001010000111101111101100",
"01111011100100111010011010000011",
"01011101100010010111100101111100",
"00011011001110110101101001001001",
"00101101010110110000000011000000",
"01011000111111110101100110000100",
"01001100001101001100101000001100",
"01000001111110111101010110000001",
"01000000101100111000101001010110",
"01010110001101000110001001101000",
"01001010110101101110010001000000",
"01010110111010001011100001101111",
"01001011001011001001011110110110",
"01100100001110100101010000000110",
"01010001110110100110011101000001",
"01101100111100101001001101100001",
"01010110001100000011010110001110",
"00011111100001100001011101001000",
"00101111100000110000001010010100",
"01101011111011001101110100011010",
"01010101101011100001111101001001",
"01001100100101001101001101111100",
"01000110000010100000010101010011",
"01010100111010011110100011011010",
"01001010001011010000100001110010",
"00101010101000001011011101010110",
"00110101000011110110110110100011",
"00110111110010000110101101100011",
"00111011101000000010101011101101",
"00110001000011001111111100101001",
"00111000001111011111110010111101",
"00000001010011001000011101000101",
"00100000011001001101001001001011",
"00110100111110111000010101000010",
"00111010001100110110110110111001",
"01110010100100110000110010110100",
"01011001000010010011000111001111",
"01100000000001010001111011000011",
"01001111101110001001101010110110",
"00011100111010100011010110101000",
"00101110001011010010010011011001",
"00000110100010010010101110011110",
"00100011000001001000000110000001",
"01010001011000110110010100110101",
"01001000011100010100011000101100",
"01111011100101001011110010110110",
"01011101100010011111101011000011",
"01001110110101010111010011001110",
"01000111001001010100101101111110",
"01101001111011001101011111101001",
"01010100101011100001110101100001",
"01011010001110111010001101101011",
"01001100110110110010101101111001",
"01101000111000011011001100011010",
"01010100001010011111100000100001",
"00001111011000111010100010000111",
"00100111011100010110100111100001",
"01100111100111101111010011100110",
"01010011100011101010010000010110",
"01001100101000000101000011001101",
"01000110000011110011111111011010",
"00001100010000010110111001001111",
"00100101110111101000011011101110",
"01100011001100101001101101101010",
"01010001010101011101010010010000",
"01100111110110111010101100010111",
"01010011101001111010111011010000",
"01100101010000001100011111010011",
"01010010010111100010011100010111",
"00100101001011100111000011101011",
"00110010010100110101001001100011",
"00111110000100000000110101111111",
"00111110110000000000100011111110",
"00111100001010011000000001000011",
"00111101110100000100111011011111",
"00001001011010001100010011110001",
"00100100011101000001101111000100",
"00101011000000101010000011100001",
"00110101001101101101111001010100",
"01011011101011111001011110001011",
"01001101100101011110101101010001",
"01110101010101011010001000001011",
"01011010011010011101101111101000",
"01110111100101110111010001011101",
"01011011100010110011101111111000",
"00110000100110011000000001100110",
"00111000000011000010110000001010",
"00011111111101100101100101100001",
"00101111101100011001001100001111",
"00101111010111111101111111000000",
"00110111011011110110011000010010",
"01100001101001100111111110001111",
"01010000100100011111110001001100",
"00100001010000101110000010100110",
"00110000010111110101101110001111",
"01100100010110110110010100000010",
"01010001111011001111110111010111",
"01010100001110011000110001000011",
"01001001110110011111001000001111",
"00000001010001111111111101101010",
"00100000011000100100010111011010",
"00000001010001011001101010101011",
"00100000011000001110101000101111",
"01011010110000101011011111100010",
"01001101000111011101111110001000",
"01010010101010110110010010011111",
"01001001000101000001110110101000",
"01111100110110100101011101100001",
"01011110001001110010110011110101",
"00101001100110000010110010110000",
"00110100100010111001000010011000",
"00111100100110000011110010001000",
"00111110000010111001011111011100",
"01010111000101011111101011001100",
"01001011010000111111001000100111",
"00010010011110011101111111001010",
"00101000111111001110101100100100",
"01001011111110111110010100010000",
"01000101101100111000111111100010",
"00111110101101001110111110110011",
"00111111000110000010111100000000",
"01011111000110100011000010011000",
"01001111010001101010110101010110",
"01011000001111010101001101011111",
"01001011110111000010011100101101",
"00100001111001111000101100011101",
"00110000101011000010011111010110",
"01000110111101011101101110101111",
"01000011001100010110010110111100",
"00111101011111100001101100110011",
"00111110011111110000110100100110",
"01000111000101011111110000001000",
"01000011010000111111001011110101",
"00000101000001011110100100101110",
"00100010001110010010011011011010",
"01111001101001111001101101110110",
"01011100100100100111100010001110",
"01010000011111101100000011111001",
"01000111111111110110000001001010",
"00110000000010001000101000001111",
"00110111101110101111010111000100",
"01010101010101110011001100000001",
"01001010011010101011011011111000",
"01000101110101000110001100000100",
"01000010101001001110000101011001",
"00100111100111111111111001101100",
"00110011100011110001101100001000",
"00000101111100001011001101100111",
"00100010101011111000011011100100",
"01100101110010101011110001100101",
"01010010101000010001011100110100",
"01010110111111111101111000101101",
"01001011001101001111100011111101",
"01100111100101110011001011110111",
"01010011100010110001110111100101",
"00000111000011011001110100001011",
"00100011001111100110011011111110",
"00111011010110110100001100101111",
"00111101011011001110101110010010",
"00111011110100001011111100111010",
"00111101101000110111011000011010",
"00001000010101011001110001110101",
"00100011111010011101100011011010",
"00111100101000001101110111011010",
"00111110000011110111111011010001",
"00010110100100110111011100011100",
"00101011000010010110001101101001",
"01011011000000010000000100010100",
"01001101001101011011101001100000",
"00111001011110110011010100111011",
"00111100011111011001011110110111",
"01000000001010111010001111001100",
"00111111110100011001111001000011",
"00010111100110010011110110011101",
"00101011100011000000110110001001",
"00010000100100010011000000001000",
"00101000000010000101001010111101",
"01010010101001011000001110010111",
"01001001000100011000110110101100",
"01100011100101010010001010101101",
"01010001100010100010101000000110",
"01001111010001100001111110111011",
"01000111011000010011010111011101",
"00110001101111111011010000101111",
"00111000100111001010010101111001",
"00111011110100100111011000001100",
"00111101101001000010000110010000",
"01110001001011011010101011011000",
"01011000010100101101101001000110",
"01111000101101011000111111011110",
"01011100000110000111001001001101",
"01111001010100001001000100111111",
"01011100011001110001000111011100",
"00111000010000111010011011100000",
"00111011110111111100110100001100",
"01111101101110110111100100001100",
"01011110100110101110100001111001",
"01110010111110000010110010110101",
"01011001001100100011101100101101",
"00001000110000100110011111011001",
"00100100000111011011111100010010",
"00101101110001000000001100011100",
"00110110100111100110010110010110",
"01001000010011110101111110110111",
"01000011111001100110100001100000",
"01001110100101101100101011011101",
"01000111000010101110110111111000",
"01010101011001000000000110001000",
"01001010011100011001100100001101",
"01001110010000000001001100011110",
"01000110110111011011111011011111",
"00110100011000011000011101000010",
"00111001111100000100100000010111",
"00101100011000111101111110110101",
"00110101111100011000011100100000",
"00110101110101110100011000010101",
"00111010101001011111111101000010",
"00111011011011110010010001001101",
"00111101011101110110110101100111",
"01100111101111110010001011100101",
"01010011100111000110101000010010",
"01110001101010000000010101010000",
"01011000100100101010011011000111",
"01000011110001001100000011000011",
"01000001100111101011001000100100",
"00100100011000000000000010111111",
"00110001111011110111011110110101",
"00001000001110110111110001101100",
"00100011110110110001010010110010",
"00011110110001011100000111010111",
"00101111000111110001100110101111",
"01011101110110110011010111111011",
"01001110101001111000001000011000",
"01001000011001110010000000111001",
"01000011111100110011111011000100",
"00110110010111101111111101110100",
"00111010111011101110111000000110",
"01101110011011000110011000000011",
"01010110111101100000000100001011",
"00011011000011001010001111010000",
"00101101001111011011111100101000",
"00011001111101000010001000100001",
"00101100101100001100011000100111",
"00111101101100101000010110111110",
"00111110100101110010101001000000",
"01001100110011000101011111111111",
"01000110001000011011101001101000",
"01010101110001101001100000101110",
"01001010100111110110111111010001",
"00101110111000000011000010010110",
"00110111001010010110011001011001",
"01000101100000011110011111011101",
"01000010100000001111001100000110",
"01001111000101110010100101101101",
"01000111010001001011011101110011",
"01100111001000111101011101110110",
"01010011010011001100110100010000",
"01000011001111010110000011101001",
"01000001010111000010111100001110",
"01000010000011110101011000100011",
"01000000101111111000111010100000",
"01101111111001100011111101001111",
"01010111101010111010110001010000",
"01110001000000010110010000000101",
"01011000001101100000000000000011",
"00001010010111101011010111011010",
"00100100111011101100011010010101",
"00111110011111010000101000101100",
"00111110111111101000001111111011",
"01000110011001010110010110001110",
"01000010111100100101010101100011",
"01011000100111101100100011111000",
"01001100000011101001000001011111",
"01110010110111101001000101101110",
"01011001001010001100100100110110",
"01110010110010010100010101000011",
"01011001001000001000000111100110",
"00001110011101100000111100001110",
"00100110111110101111101011101101",
"00101110010011011011010110111011",
"00110110111001010111101100111110",
"01011010100010000110100000101000",
"01001101000001000010001011110111",
"01110010000100100111011001111110",
"01011000110000011010001010001011",
"01111110111010000110100011101000",
"01011111001011000111101000110101",
"00001000010110011001000011001010",
"00100011111011000000000001101100",
"00010000110110000011100001010110",
"00101000001001100101110010001111",
"01011100110000111001111011100011",
"01001110000111100011110100010010",
"01010000110000001011000100000011",
"01001000000111010000110010100011",
"01000111001101110011011111001010",
"01000011010110001001001010100100",
"01001011001100000000010011100110",
"01000101010101000100011010000111",
"01101011110011010101010011010011",
"01010101101000100001111001010110",
"01100001001010110101100111101100",
"01010000010100010111000100100010",
"00001000111000101000101010100100",
"00100100001010100100100100110110",
"00111000100110011010110011010010",
"00111100000011000100000001010000",
"00110110111100011111001000011010",
"00111011001011111111101011110001",
"00110111110000101011101100111010",
"00111011100111011110000011100011",
"01111110000110111001010010101111",
"01011110110001111001001000111101",
"00000110000010010001101110000111",
"00100010101110110101100101000011",
"00011110111001101001001010110000",
"00101111001010111100101101100010",
"01000001010110001111010110011001",
"01000000011010111010110000110010",
"01001000000110000111000110101010",
"01000011110001011000110010010100",
"00001110110011001101000111111111",
"00100111001000011110101010101000",
"00110010010110100101100110011110",
"00111000111011000110110101000000",
"01010010011101110010011110000100",
"01001000111110111000100111001101",
"01001101010010011101110000101011",
"01000110011000110101001011101100",
"01111000101111111011111100101100",
"01011100000111001010100111110110",
"00101011000101011111000001111101",
"00110101010000111110101101101010",
"01000000001010000110110110011001",
"00111111110011111010010111010011",
"01101011100010010000010001110000",
"01010101100001000110111010010010",
"00111001100010111111111110001011",
"00111100100001011101110101100000",
"01101110011101100010001101010100",
"01010110111110110000010101000100",
"01000110000100010110110010011000",
"01000010110000001111001001110110",
"00111001101010100001001111101001",
"00111100100100111000101111100100",
"01100000100010001001100111010011",
"01010000000001000011101100000011",
"01000100111110011101010110000000",
"01000010001100101101001101110110",
"01000010000000111010010010110011",
"01000000101101111001001111010110",
"01110001011000001101001000101001",
"01011000011011111110011110001011",
"00100001101111010111010001100011",
"00110000100110111011100110000111",
"00010010110001000101010110110111",
"00101001000111101000011011110011",
"00111000100110000000100111110011",
"00111100000010111000000010101001",
"01101100111011010111100101001001",
"01010110001011100101100010101000",
"01111110100100011010101010001010",
"01011111000010001000110000110100",
"00011001110000110110001111011111",
"00101100100111100010010100110001",
"01110101110100000000001111101101",
"01011010101000110010110010110101",
"00110111001010110101011101011101",
"00111011010100010110111110010010",
"01010000101101010101010111111001",
"01001000000110000101100111111101",
"00101101100100101011111100100111",
"00110110100010010000110110011110",
"00110101010001101110110000001100",
"00111010011000011010100111011111",
"01010110101111100111000110000001",
"01001011000111000010000101101011",
"01001100011110010101000111010111",
"01000101111111001010001101000011",
"01110110100111111110000110100101",
"01011011000011110000111000101000",
"00011110110101101110001100101011",
"00101111001001011101100100011010",
"01011011010001100010001111010110",
"01001101011000010011100000110010",
"00101000111110100011101101000100",
"00110100001100101111011111011110",
"01110001010011100000101010110000",
"01011000011001011010101010011101",
"00101000100100000000000000000001",
"00110100000001111100001110110110",
"00100001101110011111101001110000",
"00110000100110100100101000010110",
"00011100011000111111101100101101",
"00101101111100011001010110101111",
"01101000101110000110110110011010",
"01010100000110011010010100100001",
"00001101010000101111111011100000",
"00100110010111110110110011100001",
"01010101111011111111101010111000",
"01001010101011110100001110000001",
"01010111001011101001000011101111",
"01001011010100110110010111000111",
"01010011010101000110101101111001",
"01001001011010010011000110101110",
"00001111100110100000111010100001",
"00100111100011000110110011101011",
"00110111101101110010101011000010",
"00111011100110010001111001101100",
"00011000010011100100000011111001",
"00101011111001011100100011011100",
"01010001100111011011001101010100",
"01001000100011100001001110000101",
"00101001000101111111110011101011",
"00110100010001010100000011100000",
"00111010000010111011010101011101",
"00111100101111010001111000001001",
"01100100011000100000100100001011",
"01010001111100001000110100110001",
"01100001101100000000011011011110",
"01010000100101100001101011010000",
"00100110111110010010111010100110",
"00110011001100101001011110110101",
"01100010111100111011001110010110",
"01010001001100001001111000011101",
"01111011011100110110101010111110",
"01011101011110011010000100010010",
"00011100110010010011001010010100",
"00101110001000000111101001110010",
"00011010000111110000101011110011",
"00101100110010011100011110001001",
"01001100001010001100000010110111",
"01000101110011111101100100001010",
"01001010010110111111000110111011",
"01000100111011010100100111001100",
"01001111011001011111011011111111",
"01000111011100101010001000101001",
"00100010111001110011001000111000",
"00110001001011000000011011000111",
"00010110110101010100001110010011",
"00101011001001010011100001101101",
"01000110000001011101100010100101",
"01000010101110010001101101101011",
"01000001101111100001010101100100",
"01000000100110111111101110100100",
"01110010000110110110011101101001",
"01011000110001110111010100110001",
"01101111000000000001001111101001",
"01010111001101010001001100000110",
"00110011000011000010000000010100",
"00111001001111010110011000110101",
"00011010101010110110011101101011",
"00101101000101000001111011011110",
"00010000101110100000111001011001",
"00101000000110100101001001010111",
"01001111011100000001101101000001",
"01000111011101111110110100000111",
"00000011011000111101010100000101",
"00100001011100011000000101110110",
"00011101111111010000110100111010",
"00101110101100111111100101010010",
"00100101011000000001010111111001",
"00110010011011111000001100001101",
"01011010100100100110010111110100",
"01001101000010001110001111101111",
"01110001010100010111100010110011",
"01011000011001111001000111110000",
"00110100111110100010010010011010",
"00111010001100101110111111000011",
"00010010010010011001000010110110",
"00101000111000110010100001101011",
"00001001100111111011100110101100",
"00100100100011101111110001000101",
"00000110100101111101011111101110",
"00100011000010110110100110110101",
"00111011011000011000110110100001",
"00111101011100000100101101111100",
"01000011101010110110111100001001",
"01000001100101000010001000101000",
"01101010111110011110000011111010",
"01010101001100101101011110010010",
"00011101000100011001010010000000",
"00101110010000010000110011101110",
"01101010101001001001110110110000",
"01010101000100010010100001110010",
"01001101111011011001010010010000",
"01000110101011100110001010101011",
"00011000100001001111111100111110",
"00101100000000100111100101111111",
"00000111011011011101000001000100",
"00100011011101101011110101000000",
"01101000000011001001111110000011",
"01010011101111011011110001000001",
"01100100101011011011111111110101",
"01010010000101010010000101111000",
"01010001110010011100000111111111",
"01001000101000001011001110011010",
"00110111011100101001011010000010",
"00111011011110010011010000101000",
"00000111100101001111001000101110",
"00100011100010100001001110001110",
"01101000100111110000010110010010",
"01010100000011101010101110010001",
"01111101011110000110111100100111",
"01011110011111000011000001001111",
"01001001010100110000011110010010",
"01000100011010000110111000000000",
"01011010101110100110110011111100",
"01001101000110100111100110010010",
"01101100011110001000001100010000",
"01010101111111000011101001101010",
"01111100010111110010011110100110",
"01011101111011110000001110001111",
"01110101011001011101010001100111",
"01011010011100101000111111101001",
"01111101001100101001000101101010",
"01011110010101011100111010010100",
"01001011110011110100001011100111",
"01000101101000101110000011101101",
"01111000110010011010100101101100",
"01011100001000001010100111010000",
"00011011001011111001111010100100",
"00101101010101000000100011010110",
"01110001001011110101100011100000",
"01011000010100111101111010110100",
"01010011010111000000111101100001",
"01001001011011010101100111001010",
"00001100100000010001011101010111",
"00100110000000001000101101011111",
"00100110001010010111110101111010",
"00110010110100000100110100101000",
"01100101101001011010000000010111",
"01010010100100011001101000110011",
"00010110001000001101000100000011",
"00101010110010101110011011000111",
"00101100110000010101010101101000",
"00110110000111010100111110010011",
"00100001000001110010110110111001",
"00110000001110100000011010110000",
"01011001110011000100000000001101",
"01001100101000011011000011101110",
"00010111101110110011011001100010",
"00101011100110101100110011101100",
"00111110000110001100001000111001",
"00111110110001011100000011000000",
"01000100011100001101110110111101",
"01000001111110000101000101011011",
"01100101101010001100101011110010",
"01010010100100101111110011101100",
"01010110100111011100000101110111",
"01001011000011100001100111100011",
"01001011110111101010111000000001",
"01000101101010001101010000001100",
"01001101101101010110101001110101",
"01000110100110000110001010010111",
"00111011010010111000000101101100",
"00111101011001000011111110100011",
"00011101101010000111000000000000",
"00101110100100101101010101001110",
"00000101001010000000000011111000",
"00100010010011110110001011010010",
"01000010111000000111001110011010",
"01000001001010010111111110101000",
"00000110010001110111010110010011",
"00100010111000011111011111010011",
"00000010101000000111000000011111",
"00100001000011110100110111011000",
"00001100001100110111101100101100",
"00100101110101100101101001011000",
"01100001000000011110001010001111",
"01010000001101100101100011101011",
"01101111000110001111001100110000",
"01010111010001011110000001101110",
"00001000100100101010001011010010",
"00100100000010010000000001100010",
"01010110011001111011011011110110",
"01001010111100111000111000001001",
"01101100010010111000010010011010",
"01010101111001000100000101101100",
"01010100011000011110010110111001",
"01001001111100000111101001100101",
"01001111001100010110000001100010",
"01000111010101010001011110101000",
"00000111011110110010001100111110",
"00100011011111011000111010100010",
"01000101100100010011111010011001",
"01000010100010000101100110010011",
"00100010100011010110111111000011",
"00110001000001101000110011110111",
"00010011111111000011101010010101",
"00101001101100111010111001011010",
"01101011101110101011110000010011",
"01010101100110101001101001010011",
"00001000001100110000111111011011",
"00100011110101100001101000111001",
"00101010000111010000101110011000",
"00110100110010001000001000100001",
"00011000011111000001000101111100",
"00101011111111100000011011001011",
"00101001001110100011110110010100",
"00110100010110100101101000011001",
"00000011111010010100101110100101",
"00100001101011001100111001000011",
"00110000001101110100011111011110",
"00110111110110001001110000100100",
"01100111010100101111111111001101",
"01010011011010000110100110111010",
"01001000010110100010100101100010",
"01000011111011000101001100100001",
"00010101111000000001001011010001",
"00101010101010010101101100011001",
"00111101111100001100000101000100",
"00111110101011111000101111110010",
"00010100001110001101011101100011",
"00101001110110011000011110111010",
"01100011100101010111110101000110",
"01010001100010100101001111111000",
"01111001001111000100001010110000",
"01011100010110111000100001101010",
"00110001111000010100011101100100",
"00111000101010011100111110001101",
"01101000101111010111111000111110",
"01010100000110111011110110010100",
"00111100000111001011011001001011",
"00111101110010000100101110100110",
"00111000001010001011110011110111",
"00111011110011111101011010111011",
"01101011010111011110111001011110",
"01010101011011100101101110001101",
"01001000010100000011000101110111",
"01000011111001101101110011000111",
"00011001001010101001111110000110",
"00101100010100001111111100011000",
"01011010011101101110000110001110",
"01001100111110110110011000110001",
"01010000111000101101010001001010",
"01001000001010100110010011100001",
"01101111100100100101011001111100",
"01010111100010001101110010110011",
"01000110110000100110011000101000",
"01000011000111011011111001100011",
"00100101010001001011101000000011",
"00110010011000000110101000110001",
"00111110110000111011011011011110",
"00111111000111100100011011000101",
"01001110001111011000100101100110",
"01000110110111000100011010010101",
"01101010110101011111100010011101",
"01010101001001010111111001111110",
"01100001010100010010011010100010",
"01010000011001110110010010001111",
"01100010001110011100001111111011",
"01010000110110100001001011000101",
"01010110100100001011010010110000",
"01001011000010000001100011001000",
"01101001100001000011011001111101",
"01010100100000100001011011100000",
"00001100010101101100111110010011",
"00100101111010101000000010111000",
"01101111000011001100011000101100",
"01010111001111011101011001010100",
"00010010101111100111010000010001",
"00101001000111000010001001111001",
"00010000010000000001101100111001",
"00100111110111011100001110001101",
"00011111010001000000111000001011",
"00101111011000000000100000000110",
"01111010000100010111001111011110",
"01011100110000001111011101001001",
"01011000100110100100010010011011",
"01001100000011001000010110000010",
"00110101001001000010000011011100",
"00111010010011001111101011101001",
"00111000000000100011010100100010",
"00111011101101101001001011011001",
"01101100110100110001101111111111",
"01010110001001000110001000111001",
"00011000101110011001111000100010",
"00101100000110100010001111000111",
"00110001001111100111011111010010",
"00111000010111001101000011110101",
"00011110101101000110001101100011",
"00101111000101111111001111110011",
"00000001011101110001110001100001",
"00100000011110111000010000100010",
"01101101010110110010111000011101",
"01010110011011001110000000101111",
"01010110110111010010000001011010",
"01001011001010000011110100001010",
"01101100110101010000101010111111",
"01010110001001010010001001100111",
"00110101101010110101111110010101",
"00111010100101000001101101111100",
"01110000000001111011111111100000",
"01010111101110100110101100100110",
"01000111010010111110110001001101",
"01000011011001000111101110001011",
"00000110100011100011001111011111",
"00100011000001101110101000011111",
"01011111100110100001011001011100",
"01001111100011000111000001110001",
"00001110000011100101001001110101",
"00100110101111101110000011001011",
"00101011110100101110110111100010",
"00110101101001000101000001000100",
"00011110010111011100110100111010",
"00101110111011100100100111000001",
"01011100010010111101101111011011",
"01001101111001000111001001010100",
"00010110101010001110011001111111",
"00101011000100110000100011101011",
"00111110100001011001111111010110",
"00111111000000101100100000101101",
"01101101001110011001101100110000",
"01010110010110011111101011010011",
"01101001001100110010101001011001",
"01010100010101100010101000001111",
"01001010110111000110111101101001",
"01000101001001111111100110101101",
"01011100010001100110000101011100",
"01001101111000010101101100100111",
"01111011111100011001111001101010",
"01011101101011111101110001111111",
"01011011000111001000101010100010",
"01001101010010000010111110111101",
"01111011100010100110111101100111",
"01011101100001010001110110001000",
"01110110000000110001001001001000",
"01011010101101110010110110100011",
"00110011101101101100111100111110",
"00111001100110001111100000100110",
"00110000101011101001000001000011",
"00111000000101010111101011000010",
"00101110000001010100011101101010",
"00110110101110001011011011100011",
"00100000100010011110101100111101",
"00110000000001001101110111101101",
"01001001011010000010111001100110",
"01000100011100111100110011000110",
"01011111010000111011111100111101",
"01001111010111111101101011111011",
"00111111001111100100111010100000",
"00111111010111001011100100010011",
"01001010110111110100101011000111",
"01000101001010010000111101110000",
"01001100100111101110110101011010",
"01000110000011101010000010110011",
"00010110000110110110111011111010",
"00101010110001110111101000001011",
"00110111101101000101010110000110",
"00111011100101111110111000011100",
"00000010010010100100110011101111",
"00100000111000111001001001100010",
"00000110001000110010111011011010",
"00100010110011000110001110010011",
"01111111000000000100000111010011",
"01011111001101010011001101111000",
"00001000110110001000000011001110",
"00100100001001100111100001101100",
"01100101101111010100010100110110",
"01010010100110111010011000100011",
"00001101000011101001010001001000",
"00100110001111110000110011101011",
"00110100101010110110111010110001",
"00111010000101000010001000000010",
"00000100000110110001001001110000",
"00100001110001110011111010100010",
"01101001010110100111000000100011",
"01010100011011000111100101110000",
"01001011010101000101010100110000",
"01000101011010010010010101110010",
"00000011110010100000011001001101",
"00100001101000001100111011001011",
"00100111111000000000111111111001",
"00110011101010010101101000000110",
"00111000100011011111000001100000",
"00111100000001101100101000010110",
"01101100111111010011000010100110",
"01010110001101000000010111101011",
"01110010101111000111111101100010",
"01011001000110110101010010110101",
"00010100110101000101000110111101",
"00101010001001001101101010100100",
"01101000111011101100111100010001",
"01010100001011101101010111110001",
"01001101110110010000101000000101",
"01000110101001101010110100100101",
"00010000010111101100000100100100",
"00100111111011101100110010100011",
"01011110111100011110000101011001",
"01001111001011111111010011011001",
"00000001100011111101100101000011",
"00100000100001111011000101110010",
"01000001000011010101000101101000",
"01000000001111100011010000011110",
"00001100111101110010100011000100",
"00100110001100011101110110111110",
"00100010000110011100010010000000",
"00110000110001100110011110100110",
"00001010011101010111111111001110",
"00100100111110101011000111010011",
"01101100001110101110100000000001",
"01010101110110101011110111101011",
"01100001010110000001001100100000",
"01010000011010110011000100010001",
"01010101010101001100101010010101",
"01001010011010010110010111011100",
"00111000110110011101010101011011",
"00111100001001101111101100100111",
"01110111011100111000001000011010",
"01011011011110011010110100001101",
"00001101000010010010000000011011",
"00100110001110110101110001100011",
"00111011001001000010001001001011",
"00111101010011001111101111001111",
"01111101100101101011000011110100",
"01011110100010101110001000001000",
"00001100000010010110000111101110",
"00100101101110111000100101010101",
"01000011111111001010001100011001",
"01000001101100111101001110010001",
"01100011010100111111011000101010",
"01010001011010001111000101000001",
"00011001000101111111011000110110",
"00101100010001010011110010000110",
"01111000101010000001000111001010",
"01011100000100101010110000111001",
"01100111011011110000100010011010",
"01010011011101110101111100010010",
"00000010011100100110011001011001",
"00100000111110010001101101101010",
"01000011111111000110011011111011",
"01000001101100111011111000101010",
"01101011001110010000111011100111",
"01010101010110011010100001100010",
"00101010010100100111011001010010",
"00110100111010000001110111110110",
"01111100100010100101011101011011",
"01011110000001010001000111111000",
"01011000001101100011111110001110",
"01001011110101111111111110111011",
"00011101000011101111010110110100",
"00101110001111110100111000100100",
"00010001010111101010100100011000",
"00101000011011101011111110111111",
"01000001001001010000111010011111",
"01000000010011011000111100101100",
"01101010111001111111111110111001",
"01010101001011000101001100101010",
"00100001101111010110101000111101",
"00110000100110111011010101011100",
"00100000000101101110111111111000",
"00101111110001001001001000001100",
"01101100011101111101100011111100",
"01010101111110111110010000001100",
"01100010110010101011101110100101",
"01010001001000010001011011101000",
"00101101000011100001100010111100",
"00110110001111101011101000010011",
"00001110100100011001110101111100",
"00100111000010001000011000010110",
"01101101010000000011101101110011",
"01010110010111011101011000100111",
"00011001010010010000000010111101",
"00101100011000101101011100111100",
"01101111111010011011000010011100",
"01010111101011001111001110100100",
"01000010100101010000011000001000",
"01000001000010100001110011000001",
"01010010001000101101011000011001",
"01001000110011000010101111110111",
"01100111010111010011001010110110",
"01010011011011011111011010110010",
"01001111100111100010011000100011",
"01000111100011100100011100110011",
"00001101010001101111100001100100",
"00100110011000011011000011011111",
"01100100111100111110001110101010",
"01010010001100001010111110001000",
"01011011101001111000100000010001",
"01001101100100100111000000010100",
"01010001010000111001101101111101",
"01001000010111111100011010001000",
"01001000010001111101100111010100",
"01000011111000100011000010010110",
"01110100101111110111111001000111",
"01011010000111001000111101110010",
"01001001111010111010110101001000",
"01000100101011011010111101111001",
"00101111101101101110001001101111",
"00110111100110010000000000101110",
"01110111001100011110010010100000",
"01011011010101010110011100001010",
"00001101111010000001010001000011",
"00100110101011000101101011001011",
"00011010111011111111000101010110",
"00101101001011110100000000010011",
"00100001100001000101101011110010",
"00110000100000100010100011001111",
"00001010011100100110101110011110",
"00100100111110010001111000011111",
"01110011001001100011000011100100",
"01011001010011100100001110011101",
"00111110100100110101000010100110",
"00111111000010010101000101111101",
"00011011110100010001010010110111",
"00101101101000111001011110001111",
"00110100010010110011111110000011",
"00111001111001000001101010101010",
"00101001011110110101000001100000",
"00110100011111011010010101101010",
"00111101100011100111111011110100",
"00111110100001110000110110111001",
"01010100011000100010111101111100",
"01001001111100001010000110100100",
"00010101111100110010100101011100",
"00101010101100000110110000000000",
"00100000010110010011101010011001",
"00101111111010111101000110101000",
"00000001011100000100100000111000",
"00100000011110000000010000111101",
"00100100100001001100011011011001",
"00110010000000100101110111010010",
"00001101100110010111011000001100",
"00100110100011000010011101010000",
"00011010101110010100100011110110",
"00101101000110100000000001100110",
"00010100011011100111011101110101",
"00101001111101110001001111101100",
"01010000001011100111110000010100",
"01000111110100110101100100100101",
"01101100110111000001111100001111",
"01010110001001111101101100001110",
"01111011110010111010101000101100",
"01011101101000010111010110010000",
"00011111110011001010001000110111",
"00101111101000011101011111000100",
"01111010001000110001011101110011",
"01011100110011000101010011101011",
"01100000101111111000110111010110",
"01010000000111001001010111001101",
"01111011011101000010101001001000",
"01011101011110100000001100110110",
"01001011011001101011001011110000",
"01000101011100110000010100111011",
"00101001000001110110011110101011",
"00110100001110100010111010001011",
"01110000001100111010100010001111",
"01010111110101100111010101110000",
"00010101010100100110000000111000",
"00101010011010000001000111000101",
"01011000101111100100101000011010",
"01001100000111000001000101000100",
"01100111011001011000110100101111",
"01010011011100100110101001010000",
"00100011001110100111010001111011",
"00110001010110100111101001000110",
"01110011101011100011101101110000",
"01011001100101010101011001101100",
"00001000111010011110100000100001",
"00100100001011010000100000101110",
"00101101101011001110000000011010",
"00110110100101001100000101000111",
"01100110110101000110110001010101",
"01010011001001001110010011110111",
"01000111011111010011100011000111",
"01000011011111101001101101101011",
"01001001011111011111010011010001",
"01000100011111101111100111100010",
"00011011000111111010101111011000",
"00101101010010100010110110000000",
"01110000111110001000100100100111",
"01011000001100100101110001011101",
"00000111000011000111001111000101",
"00100011001111011001111010111100",
"01101111100000011101101101010100",
"01010111100000001110110011001111",
"00000110111010111011001010000100",
"00100011001011011011000101100111",
"00100111011001011010111001011110",
"00110011011100100111101111010101",
"01110000111100100010001110001101",
"01011000001100000000110011101100",
"00101011011100000111100101011101",
"00110101011110000001110110011001",
"00110100111111110010010001101010",
"00111010001101001011011100111111",
"00001011101010110110110010000011",
"00100101100101000010000100010001",
"00111111110111101111000011010010",
"00111111101010001110110101011110",
"00000101001011011010000001111110",
"00100010010100101101001111111110",
"01111000100001111000101110010010",
"01011100000000111011011111110101",
"00111011101010101001101011111110",
"00111101100100111100011001101111",
"00100100111110100100001010110101",
"00110010001100101111101010000111",
"01110010101010101010001100000101",
"01011001000100111100100111101001",
"00011100011010100010100011010101",
"00101101111101001101011000011001",
"00100000011011100110110011111101",
"00101111111101110000111010000000",
"00111110000100010101010111110101",
"00111110110000001110001101110001",
"01000101011100011001000010000000",
"01000010011110001010110101110000",
"00010000101000100001010110001100",
"00101000000100000000100110010011",
"01010011011000111011011000101110",
"01001001011100010111000100011101",
"00011110001011111101101010011010",
"00101110110101000010110100000101",
"01111000000001111010001010111011",
"01011011101110100101011100100001",
"01110110100111100010101010101001",
"01011011000011100100100100111100",
"00010001110111100001011000001010",
"00101000101010001001101001100110",
"00000000111100011000101011011100",
"00100000001011111101010101100001",
"00100100010010110000101011000011",
"00110001111000111111110100001110",
"01111000101100101000001001011111",
"01011100000101110010100011010010",
"01001000011011101100001110100011",
"01000011111101110011101101100000",
"01101101110010001111111110010100",
"01010110101000000110011000011010",
"00010011110100100010111000111000",
"00101001101001000000010110001100",
"00111001011001110100110011001011",
"00111100011100110101011000110111",
"01110100110101010111001101011001",
"01011010001001010100101011101101",
"00000011010101000000100110001100",
"00100001011010001111101111100111",
"01000000010100101111111101001111",
"00111111111010000110100101110101",
"00011100001110110010000110110111",
"00101101110110101101111110101101",
"01110100010001100010110100011001",
"01011001111000010011110101110110",
"01101011110000110111100010101100",
"01010101100111100010110110011100",
"01010001001110100100011000100001",
"01001000010110100101111100011100",
"00101011101000100110100101111110",
"00110101100100000010111011011010",
"01010110011001111110011010011111",
"01001010111100111010011100010011",
"01111000011110010010010100101110",
"01011011111111001000110010100010",
"01100111010011010000010001111101",
"01010011011001010001100001001100",
"01111011011000100010100101010100",
"01011101011100001001111001011110",
"01101011001000111100100000110011",
"01010101010011001100001110000110",
"00000011101101110010110101010010",
"00100001100110010001111101111110",
"00011011110100001001011001010001",
"00101101101000110110011000010101",
"00101001001101010001111000101001",
"00110100010101110101001111111001",
"01001001001010001011110111010010",
"01000100010011111101011101000010",
"00101100011100101010101111011101",
"00110101111110010011111100100000",
"01111100100110001101010001010111",
"01011110000010111101110101100101",
"01100111010110001001100001101100",
"01010011011010110111100110010010",
"00100100011110100100111010011000",
"00110001111111010010001100110010",
"01110011001101101111111100000000",
"01011001010110000111000100010010",
"01111001001101101010111001110110",
"01011100010110000100000101101011",
"00100101011010111101100101110100",
"00110010011101011011011111011110",
"00010111100000100000100111000100",
"00101011100000010000001111011010",
"01110001111010010011000011010110",
"01011000101011001100010001010110",
"01101101110110101001110100011000",
"01010110101001110100011110100100",
"00000101010010110000100101011000",
"00100010011000111111110001000010",
"00000101101110110101111100001110",
"00100010100110101101110110111100",
"00100111010000011110100111100011",
"00110011010111101100110111111000",
"01111010001000000111110010110010",
"01011100110010101011000110010000",
"00001001000011110110100010011010",
"00100100001111111001101011110110",
"01100111100101001110100100110010",
"01010011100010100000111101100100",
"00010110010110111001111001101001",
"00101010111011010001110011010110",
"01111101010101011001010110110100",
"01011110011010011101010100100111",
"01010011010110000110000111011110",
"01001001011010110101101111100111",
"01100111100101011110010010001011",
"01010011100010101000001110110111",
"01111101010001110010111101010000",
"01011110011000011101000000000100",
"01111110111110101100101101011100",
"01011111001100110010101101011110",
"00111101111111011100101100101010",
"00111110101101000011110011010000",
"01110101110000000101010001111111",
"01011010100111001110011011101011",
"01100110010001111100111111011001",
"01010010111000100010101011110000",
"00111001010111111111010001111111",
"00111100011011110111000100101010",
"01100000111001000001110010110010",
"01010000001010101110000000001111",
"01101001111111101111110100101011",
"01010100101101001010100101011000",
"01010101001100001000101011010000",
"01001010010101001001011100111000",
"00001010000110010011101011011011",
"00100100110001100000111011000110",
"00110011001001111011101011111101",
"00111001010011110011011110011100",
"00000001101000110011011010101110",
"00100000100100001000100111010010",
"00000110101100100000111100110010",
"00100011000101101111100000000111",
"00011010100000000101001101101001",
"00101101000000000010100110101101",
"00100110000111011000010101000110",
"00110010110010001100111111000000",
"01111001111010010000111000110011",
"01011100101011001011011110000000",
"00010011101101110000000111100000",
"00101001100110010000110101010100",
"01001011100010010101111010111011",
"01000101100001001001101000101111",
"00010001011010110001011111110111",
"00101000011101010101001011111110",
"00000101101000000011001010110110",
"00100010100011110011001001101000",
"00111001011000111111101111010011",
"00111100011100011001011000000111",
"00010110101101100010000101001111",
"00101011000110001010111101010000",
"00001011010110111001000111000100",
"00100101011011010001011000000010",
"01100000101001011110010110110110",
"01010000000100011011100011001001",
"00010000110101101001111000000001",
"00101000001001011011111001101000",
"00010100011010101111101001011110",
"00101001111101010100001110001100",
"01001000001110101100111011101000",
"01000011110110101010111100111010",
"00100111001100100011110001101011",
"00110011010101011001101110101100",
"00010001110000001001000000010010",
"00101000100111001111111100110110",
"00011011100100110011000011000110",
"00101101100010010100001010100010",
"00001110110010000010000011110110",
"00100111001000000000110100101110",
"00001111000001111011111101100011",
"00100111001110100110101011010000",
"00011010100011011111110000100010",
"00101101000001101100111110101100",
"01001100110001011110110000100000",
"01000110000111110010101010110001",
"00000100110010000001001111100010",
"00100010001000000000011111110011",
"00000000110101011100101111111100",
"00100000001001010110110100111011",
"00000110001001011110000010011111",
"00100010110011100001000111000111",
"01100101101011000011000010010100",
"01010010100101000111010110101111",
"01101010110101001100100100100111",
"01010101001001010000100011111010",
"01011011010101100110101101110000",
"01001101011010100100101000001001",
"01101111110001010110101101110000",
"01010111100111101111011011101010",
"00011101111111001000010000100101",
"00101110101100111100100010001100",
"01011100111110011010001000011110",
"01001110001100101100000100010001",
"01110110011101110111101010100010",
"01011010111110111011010000010101",
"00111000011111001101011110001110",
"00111011111111100110101010000101",
"00000011000101110010011101100100",
"00100001010001001011011000100001",
"01110000011000001000100011010101",
"01010111111011111100000001101000",
"01001100001100111101100101101110",
"01000101110101101001001010011010",
"01001110101000001000011000011111",
"01000111000011110101011110101010",
"00000001110010111010000011001100",
"00100000101000010111000111011000",
"01010001110101000000110000100100",
"01001000101001001011111110011101",
"00001000000001001000000111110010",
"00100011101110000010110111011001",
"00011000100000011100001000011100",
"00101100000000001110000001001001",
"01011101001011111001110111101000",
"01001110010101000000100001100101",
"01101000101010100110011110101000",
"01010100000100111011000000110010",
"00101001010110000110000000011101",
"00110100011010110101101011110011",
"01110001100110101001100001000111",
"01011000100011001010101110011010",
"00110000111001010011011010010000",
"00111000001010110100100110000001",
"01010000100010101001110010001000",
"01001000000001010011001100111001",
"00000011010110110010100001011001",
"00100001011011001101110100010001",
"01001100011110000110011101010110",
"01000101111111000010110001011000",
"01011111010100101011110101111110",
"01001111011010000100010100110001",
"00010010011000101110011110111100",
"00101000111100010000001110010010",
"01100111000001100110001101111001",
"01010011001110010111101101010010",
"00101100000110001010100110011111",
"00110101110001011011000011010010",
"00010111001010101111101110011110",
"00101011010100010011011101111000",
"01100111110111000010111101110101",
"01010011101001111110000101001101",
"00110010001111101000101000111110",
"00111000110111001101101110100011",
"01111100110101110010110000110011",
"01011110001001011111010101000111",
"01010010101100001111100010011100",
"01001001000101101000000110111111",
"00001101100101001111010110101110",
"00100110100010100001010100101101",
"01101100100111001001011110100011",
"01010110000011011001001110000000",
"01110000101011010111110011000001",
"01011000000101010000010010011101",
"01101010100011101001011111001100",
"01010101000001110001100101111110",
"01100011000101000001001001000101",
"01010001010000101011001000000000",
"00101001001010100101010001010000",
"00110100010100001101000100000010",
"01101101101001011011111100110001",
"01010110100100011010011111011110",
"01010011011101001001101100011011",
"01001001011110100011110011110011",
"01110101010111100010110110111110",
"01011010011011100111110110010011",
"00111100010001100100010101010000",
"00111101111000010100101100111000",
"01010101010000000011101111100111",
"01001010010111011101011001101010",
"01000111001100100011100111100011",
"01000011010101011001101000100111",
"01000100010010101100011101000011",
"01000001111000111101011100100110",
"01101101110000011111111000000011",
"01010110100111011001010000011101",
"00100100011000011101011111001011",
"00110001111100000111001011111010",
"00101100111101010010111011101011",
"00110110001100010010011101011101",
"00010111000110100101111000100001",
"00101011010001101100101010101011",
"00010101111111000111000000010010",
"00101010101100111100000101100110",
"01011101110110100110010101111100",
"01001110101001110011001001011011",
"01100111101001001111101010101001",
"01010011100100010101000101101010",
"00011001010101111001100001101100",
"00101100011010101110111001000000",
"00101010010100101100110011010010",
"00110100111010000100110110100100",
"01000110111101111011100000101000",
"01000011001100100001000101001111",
"00101011101110101000000000101000",
"00110101100110101000000110000011",
"00010001010110010011000001001011",
"00101000011010111100110000010000",
"01110011000100000110000111000111",
"01011001010000000100000100100011",
"01000010111001010111101111000111",
"01000001001010110110001101011011",
"01111001001101010101111111000000",
"01011100010101110111101011110010",
"00100101010011101110110000000101",
"00110010011001100010100000010001",
"00111111101111001010011111111010",
"00111111100110110110010101101110",
"01001011111001100101100001011101",
"01000101101010111011010110100110",
"00110010111000111110000110110100",
"00111001001010101100100111110101",
"00101100010110010011111110011101",
"00110101111010111101010001100001",
"00111100100100111101010100011110",
"00111110000010011000111100101101",
"00011101011100100111100110000000",
"00101110011110010010010101000010",
"00001111011011010101000111100010",
"00100111011101100111101110100110",
"01100101101111100010100101101110",
"01010010100111000000001111011110",
"00001011000110000011100010110001",
"00100101010001010110011110100111",
"01100010111000011110110011111101",
"01010001001010100000110111101011",
"01011011000111000101011100101101",
"01001101010010000000111011010100",
"01000111010111100111111000000010",
"01000011011011101010100010100100",
"00111000001000100010100011100101",
"00111011110010111011111101000011",
"00100010010011101001000100010000",
"00110000111001011111010101110101",
"00001011101010010100010101000101",
"00100101100100110011001000100110",
"00100101111001000010011011101000",
"00110010101010101110001111100001",
"01000110101100000110100011011011",
"01000011000101100100010010010001",
"00111000100111100111010000110000",
"00111100000011100110101001001011",
"00111100111111101000010100001001",
"00111110001101000111111011000100",
"01011100101011001101100011101110",
"01001110000101001011111000110001",
"00010110011110001101100110101100",
"00101010111111000110011001011011",
"00100100101000110111111110110011",
"00110010000100001010101000100100",
"01110110000001000111000101011010",
"01011010101110000010001001010001",
"01000000110010111010011001111111",
"01000000001000010111010000011011",
"01101011100110110011011111011011",
"01010101100011001111010000100001",
"00100001101111101111000110000010",
"00110000100111000101010111011100",
"01010010001001001101011011001010",
"01001000110011010110110001100110",
"01011110101010111001100110100010",
"01001111000101000011010010001111",
"01100100101001000110110101001001",
"01010010000100010001001100011001",
"01001011010110100011011010001011",
"01000101011011000101101001000010",
"00000011111110101000010110100111",
"00100001101100110001001001110101",
"00100100011000010001010101000011",
"00110001111100000000101101010110",
"00010111010000001000111011101000",
"00101011010111100000011001001000",
"00110110110111100110011101011011",
"00111011001010001011100101000010",
"01010000101110100101010011100000",
"01001000000110100110111110010100",
"01010011110101000110010000000110",
"01001001101001001110000110111101",
"01010100010100001110000011011100",
"01001001111001110011110111110010",
"01100000001001111010011011000011",
"01001111110011110010101100011110",
"00111001100100101000110101110101",
"00111100100010001111011001100110",
"01011111011010010001100110001101",
"01001111011101000100100000011101",
"01000011000010011001001111000000",
"01000001001110111010101101010011",
"00010100101011101110010010100010",
"00101010000101011001111011011101",
"00100110110001111001011110001111",
"00110011000111111101011000110010",
"01111011001010111011110010100101",
"01011101010100011010110101101111",
"00110110111111010111010110110010",
"00111011001101000001111001110101",
"00110010011100001101110011010100",
"00111000111110000101000011100010",
"00100001000011111110001110001110",
"00110000001111111110110100000111",
"01111101101011011101111010001101",
"01011110100101010010111010011001",
"01101011000011110101000100000101",
"01010101001111111000101100110100",
"01011110000011100110100010010111",
"01001110101111101110111110100011",
"01011010010110101011011101111011",
"01001100111011001010000000001011",
"00000001100010000010101010110001",
"00100000100001000000010100101110",
"00000010101100011110100001001010",
"00100001000101101110011110000111",
"01010000010111110010100011010101",
"01000111111011110000010000110001",
"01000010010100111101000100110000",
"01000000111010001101110011101110",
"01101110010011010010000000100101",
"01010110111001010010011111000000",
"01110010000111100001101001011000",
"01011000110010010010111010101111",
"00010100011110001010011111111011",
"00101001111111000100110100100110",
"01001100111110001011100111000111",
"01000110001100100110110111001110",
"01010110110000101000011110100001",
"01001011000111011100101111110111",
"01011111110100101101111010000110",
"01001111101001000100101001001000",
"01010000111100110011111101101111",
"01001000001100000111010000000010",
"01111011001000111001110011100101",
"01011101010011001010100001110010",
"01110111000100110110110101101110",
"01011011010000100100010110000011",
"00000111110100011010011011001010",
"00100011101000111101000010101100",
"01001011110111011111000111000101",
"01000101101010001000110010100010",
"01001010111001111101000101110100",
"01000101001011000100000111111010",
"01011100001000101000011110100110",
"01001101110010111111101011000010",
"00101100000001011001100010001000",
"00110101101110001110111100010010",
"00000100011110100101111011101001",
"00100001111111010010101101110010",
"00111011100010111010000100110100",
"00111101100001011011000000111110",
"01101111000011110010110001001001",
"01010111001111110111001010100110",
"00011001001010010100001110001011",
"00101100010100000010100110001100",
"01100010010100110011100011000011",
"01010000111010001000100100010110",
"01101010001110101110100011101110",
"01010100110110101011111001110101",
"01010000001001101011100100111101",
"01000111110011101001100000101001",
"00010100110001000001010110011000",
"00101010000111100110110100001110",
"00001011010010101100110001111100",
"00100101011000111101101000010100",
"01001101110101001001011111001011",
"01000110101001001111010111010101",
"01101001010110010011010100010100",
"01010100011010111100111010101010",
"00101000001011110100111101000110",
"00110011110100111101100011100111",
"00000001010110111001000101001110",
"00100000011011010001010111000010",
"01101100000010110001110101011110",
"01010101101111001011011100001101",
"01111000100011100111100000011100",
"01011100000001110000101001111010",
"01000011101011110110001001111111",
"01000001100101011101010010101010",
"01011010010110000011110110000100",
"01001100111010110100100000100001",
"01101010101011001001001001110100",
"01010101000101001001111111011011",
"01011000001010000000101001111010",
"01001011110011110110100010110001",
"00100111010100001111011101001011",
"00110011011001110100101001011101",
"01000001011011110001101000010101",
"01000000011101110110100000011101",
"00110111111110101110100100000000",
"00111011101100110011010111110100",
"01111000010001000011011010111010",
"01011011111000000001111101000010",
"00111100100100101011011011111010",
"00111110000010010000100111001100",
"00101111000011100101011001101110",
"00110111001111101110001101110101",
"00001000011100001010100011000000",
"00100011111110000011011000001010",
"01111001111101100010011111100010",
"01011100101100011000000100110111",
"01011100001110000110010100101011",
"01001101110110010100010001111010",
"00110100011101100100000101001000",
"00111001111110110001010010001001",
"01111110011100001000011011001100",
"01011110111110000010010010000111",
"00010111110001000000011001011111",
"00101011100111100110011011100111",
"00100011100001010110110110010001",
"00110001100000101010111110010010",
"00010111100110011100101001010111",
"00101011100011000100110111001000",
"01111010000101110011111100100011",
"01011100110001001100010110010101",
"00001101110000000101011010000000",
"00100110100111001110011110111100",
"01100111110000001000001110010101",
"01010011100111001111101000011110",
"00001110110110110101010010111011",
"00100111001001111000110111010111",
"00011001000010110010001011111100",
"00101100001111001011101011011011",
"00110101100101010001101101100000",
"00111010100010100010011010100101",
"00001110101011101011101101011000",
"00100111000101011000110100110011",
"00000010011001000101100000010000",
"00100000111100011100011011100001",
"01011101110001000110101010100110",
"01001110100111101000111101100110",
"00010000000010100100110010100110",
"00100111101111000010100101000101",
"01101110011011110111010101101111",
"01010110111101111001011101011100",
"01010110010100101110001011000010",
"01001010111010000101100110111010",
"01010011101110011010111100100101",
"01001001100110100010101011010111",
"01001000110001111011001011110011",
"01000100000111111110000100101010",
"01000000111111110111010100110110",
"01000000001101001101001111011001",
"00101011111000011011100110011111",
"00110101101010011111101010010101",
"01110000000110001010101000111110",
"01010111110001011011000100111001",
"00000010011011101000111101001100",
"00100000111101110010000001000110",
"01100011110111001010001010011111",
"01010001101010000000110100101111",
"01101000010111001110000011111001",
"01010011111011011100101010110111",
"00111111000000010100011001000110",
"00111111001101011110101100010110",
"00010010111010101111100100001101",
"00101001001011010110110100000011",
"01101000011100101011111001111110",
"01010011111110010100100010110001",
"01000111011100011110111100000110",
"01000011011110001101111000010010",
"00001100111000010010000011110000",
"00100110001010011100000100001111",
"01000100101010110010001110101001",
"01000010000101000000000110010100",
"01111011111010000011000001001111",
"01011101101011000110010100110100",
"00001011010100011010011110111100",
"00100101011001111010101111101101",
"01011100011011110010101000001001",
"01001101111101110111000001011110",
"00011111011011011001110111100000",
"00101111011101101010001100011010",
"00100010111010110111001000010011",
"00110001001011011001100110101000",
"01010110100001100110100100101100",
"01001011000000110010101010001111",
"00101101001011011111010001100000",
"00110110010100110000011011100110",
"00001010101010111111010110101000",
"00100101000101000101110001000110",
"01100101011000011011110111100111",
"01010010011100000110010100110010",
"01000110001110010001011101011101",
"01000010110110011010110101011100",
"01000000010000010001000100001000",
"00111111110111100101000101000001",
"01110100000100000111100100111111",
"01011001110000000101000011000011",
"01001000100111010110111101101101",
"01000100000011011111010011101011",
"00011110000001010111101110101111",
"00101110101110001101101100011000",
"00000100000110101100010111100101",
"00100001110001110000110101110000",
"00110111000011001110010011011100",
"00111011001111011110101100000100",
"01110100010110000101111001110001",
"01011001111010110101101000001010",
"01010111110101000111010100001011",
"01001011101001001110100001011000",
"00110101010101111101001110101000",
"00111010011010110000111010000011",
"00000011101101100010111010101010",
"00100001100110001011010011101001",
"01101111111011010100001000001110",
"01010111101011100100010001100001",
"00110111110001100110001011110100",
"00111011100111110101101001110001",
"01100111100100101101000101001010",
"01010011100010010001011000010101",
"01011000010010100010001100000111",
"01001011111000110111101011001111",
"01110110110001111010100100111010",
"01011011000111111101110101000110",
"01111010011111011100101001010111",
"01011100111111101110010010001110",
"01000000101111001110000110000101",
"01000000000110110111110100100000",
"00111110001110011001100001000001",
"00111110110110011111100100011010",
"00000111010111101110101101000111",
"00100011011011101110001100110111",
"00000101011010000000010100101110",
"00100010011100111011011100100001",
"00111010001000011100100010010000",
"00111100110010111000001010110101",
"00010010101100001001001100000011",
"00101001000101100101011010000101",
"01100001110101110010111100110111",
"01010000101001011111011001110001",
"01011001100011110110011001110000",
"01001100100001110111101100111110",
"00110101100111000000010100010111",
"00111010100011010101000100110001",
"00111000010111011001100001100011",
"00111011111011100010110101011101",
"00000110101111010101101011010001",
"00100011000110111010111100000101",
"01000000010001111111101010111111",
"00111111111000100100001100110110",
"00011101101111110101011001001010",
"00101110100111000111111100010111",
"01001100111101100111001000101110",
"01000110001100011001101111111111",
"00000000100010010000101111001000",
"00100000000001000111001000011111",
"00010001110011111100111110001001",
"00101000101000110001100000100110",
"00010101100100111110000110011011",
"00101010100010011001010011111101",
"00011110100011101000011101110111",
"00101111000001110001000111000001",
"00010101111010101001010101101111",
"00101010101011010100100000111100",
"01001100101000001100011001111000",
"01000110000011110111010001100010",
"00010010111001101110010111101000",
"00101001001010111110101001100000",
"01101101101111110000101001111010",
"01010110100111000110000000010011",
"01001100011101010101111001000111",
"01000101111110101010000010110100",
"01001000001111101011100110010000",
"01000011110111001111011100001110",
"01110001011101010011100100100100",
"01011000011110101000110110111100",
"00111100011000101010000001010101",
"00111101111100001101110110100100",
"01011001000010000000101001101110",
"01001100001110101001111001001110",
"00010100101011001100001101011100",
"00101010000101001011010011101000",
"01110110110011001100010110111111",
"01011011001000011110010111010000",
"01010011100001011101010011000110",
"01001001100000101110001000010010",
"01010101011010011010010011100001",
"01001010011101001001000100010011",
"00110101000001100101111000000000",
"00111010001110010111011110001100",
"01011010111001001100000000001101",
"01001101001010110001110100110011",
"01011010110100011010101000010000",
"01001101001000111101000111110011",
"01101111001010000010011010010000",
"01010111010011110111101000000101",
"01101101100101010101001100010001",
"01010110100010100100000001101110",
"00111100101010001101100101000111",
"00111110000100110000001100101010",
"01001000101101111000110100000000",
"01000100000110010100011101110110",
"00100011001100010101100000101000",
"00110001010101010001001010111000",
"01110101000001100111000110101011",
"01011010001110011000010100011110",
"01001111011101001110011111010001",
"01000111011110100110010000101101",
"01100011011110010101001011100111",
"01010001011111001010001111001101",
"00010010110001011100011111110101",
"00101001000111110001110000100101",
"00011100011010110101100111111111",
"00101101111101010111010101101111",
"01100100000000100101111010101111",
"01010001101101101010111111111001",
"00100100100101011001011101111111",
"00110010000010100110000000011001",
"00110001111111110011101110011011",
"00111000101101001011111101110101",
"00000010100100001110011000100110",
"00100001000010000011000000001000",
"00111010100000000010110011101110",
"00111101000000000001011001110100",
"01111110101000000000001000010011",
"01011111000011110001110010101010",
"00010101011101111100110000001111",
"00101010011110111101110101111010",
"00101000001111110011011101101000",
"00110011110111010011111111101000",
"01001011000101010110000001011010",
"01000101010000111000110100101000",
"01011101101101101000010110011111",
"01001110100110001101100101010110",
"00011001101101000111000010001100",
"00101100100101111111100101111101",
"00000111011110000000000010110000",
"00100011011110111111100000111000",
"01011101101110111010001000100100",
"01001110100110101111100101110011",
"01110010101111000111101011111011",
"01011001000110110101001011100101",
"00011100001001001100010000001100",
"00101101110011010110000010111000",
"01010100100010000110011111100011",
"01001010000001000010001011010101",
"01000110010000100100111111000001",
"01000010110111110000100001110111",
"01110001100011100110100011101110",
"01011000100001110000001101001000",
"00001001100011101100010111100011",
"00100100100001110010111101010010",
"00100001001001110000111111001110",
"00110000010011101100110111000011",
"01001100011000000001001011111110",
"01000101111011111000000101110110",
"01111000101101101110110001110011",
"01011100000110010000010001011110",
"00001110101111000110001011011111",
"00100111000110110100100011110101",
"00001001000010001110110001000101",
"00100100001110110011100011110110",
"01000001011011100111100101110011",
"01000000011101110001010011110101",
"00110001111011011011101100000111",
"00111000101011100111000011001000",
"01111110000011110101110111110000",
"01011110101111111001001111010111",
"00010000111000110110000101000101",
"00101000001010101001100111001101",
"00010101011001110000110111101111",
"00101010011100110011010100100011",
"00010000110101010010010111100110",
"00101000001001010010110011101101",
"00101101010011101011101101000100",
"00110110011001100000110011110010",
"01111001011010010110110010011110",
"01011100011101000111001110011111",
"00110101011010101011110101100101",
"00111010011101010010001110111000",
"01011111010011011111011011011111",
"01001111011001011001111110010001",
"01111011111110100101001011000101",
"01011101101100110000000001000101",
"01101111111010101110101001010011",
"01010111101011010110011110010100",
"01011101111011011111100011110010",
"01001110101011101000011101111110",
"00010001011100100001111011010100",
"00101000011110001111011010100111",
"00011000001010100010000110111011",
"00101011110100001011000111111111",
"00101001000000110101100101001101",
"00110100001101110101111100111101",
"01101111001010001010010001110011",
"01010111010011111100011110100001",
"00110001110111101001001001000111",
"00111000101010001100100110001001",
"00110000011110110101100111111101",
"00110111111111011010101001000100",
"01001100111001000100011010010111",
"01000110001010101110111110111111",
"00100100100110110000110101000010",
"00110010000011001110000011001001",
"01001100101000000001111000001001",
"01000110000011110010100100101011",
"00100001011011001010111001111010",
"00110000011101100010011010111100",
"01101010110111010101110100000011",
"01010101001010000101010000011100",
"00111110001011101000011011110111",
"00111110110100110101111110111101",
"00101010111110110111010001011101",
"00110101001100110110011110110010",
"00001100000001000110110011010010",
"00100101101110000001111100101011",
"00001010100011101001100111110101",
"00100101000001110001101010000100",
"00100011101100100110000011010000",
"00110001100101110001101010011100",
"00011010110000001100111110110001",
"00101101000111010001100100100011",
"00010011100101111000011000111011",
"00101001100010110100010000101110",
"01100101001000001101101001000100",
"01010010010010101110110010011101",
"01001100101011101000101010111001",
"01000110000101010111100001100011",
"00010001101001101110010000101011",
"00101000100100100010100001100001",
"01110110000001000011101110001001",
"01011010101101111111110011100101",
"01100010000101011001100010101000",
"01010000110000111011000111111111",
"00100010011111000000101000010001",
"00110000111111100000001100001110",
"00100011010100101111011011001101",
"00110001011010000110010011000101",
"01011011011111110000010101000110",
"01001101011111111000001010000100",
"01010111111001101100011101110110",
"01001011101010111101111100001010",
"00000010101000001110110110101101",
"00100001000011111000010111100000",
"01010111011110010101100000001011",
"01001011011111001010011001101000",
"01000111110100011011000111001001",
"01000011101000111101010011110111",
"01100000100011101110011010011111",
"01010000000001110011111011001111",
"01101000111010110111011011011111",
"01010100001011011001101101101100",
"01011111111110111101001110000100",
"01001111101100111000100110100001",
"00001001100100100011111111101100",
"00100100100010001101001000100110",
"01011000000101000001101101010011",
"01001011110000101011011111110100",
"00010001110110100110010111001100",
"00101000101001110011001001111001",
"00111010000011011001100111101001",
"00111100101111100110010011100011",
"00100100111110000110000111101010",
"00110010001100100100111001000111",
"00110110011101010111001100001110",
"00111010111110101010101101010000",
"00000110101011011011011111110011",
"00100011000101010001111000001000",
"01000110011001010001000001100101",
"01000010111100100010100001100100",
"00100001010100101101000000010010",
"00110000011010000100111101101110",
"01000100110111000011111011101010",
"01000010001001111110011100110001",
"01110001011000001000010011000010",
"01011000011011111011111000111100",
"00101101010101110011110011100100",
"00110110011010101011110001011100",
"01001111011010101101100011100000",
"01000111011101010011001000010001",
"00010101000100101110010110010011",
"00101010010000011110101111101011",
"01001000000110000000110010010101",
"01000011110001010100101100001010",
"01100011000000100101111100011011",
"01010001001101101011000001000101",
"01111010001100111011111111010111",
"01011100110101101000001101010101",
"00010100110001101001011101001110",
"00101010000111110110111101110111",
"01110100101010010100001101000110",
"01011010000100110011000101001000",
"01110000001101111111101101100000",
"01010111110110010000011000011110",
"01110110110111000010111111110110",
"01011011001001111110000101111110",
"00010111001001010100110101011000",
"00101011010011011011011000110111",
"00010011100010101111001000101101",
"00101001100001010101110001011001",
"01010010010110110011010100111101",
"01001000111011001110010000001001",
"01101111000011000001010011001110",
"01010111001111010101111010010110",
"00010110001010111101111111011010",
"00101010110100011100001011101011",
"00101001110101001000110101001000",
"00110100101001001111000111000001",
"00110110110111011100011010011000",
"00111011001010000111110000111011",
"01110110101110101100011001111010",
"01011011000110101001111010100001",
"00010010110000000000010000101000",
"00101001000111001100011000100010",
"00010110110110011001101000011100",
"00101011001001101110010001110000",
"01101010110101000001111101111011",
"01010101001001001100011100100000",
"00101000101100111111111111101000",
"00110100000101111100101000000110",
"00111010010110101010000001010000",
"00111100111011001001001110000011",
"00001111110011001000000101100101",
"00100111101000011100101011001001",
"01011111001010010111001011110111",
"01001111010100000100011010110010",
"01000001000010000101100001000011",
"01000000001110101101001110101010",
"01010110001100011001000111001010",
"01001010110101010011010101010100",
"00000101111001001001011100101101",
"00100010101010110000110111101000",
"01000111100100100001011010001101",
"01000011100010001011111011001011",
"00101101110100110111111111101101",
"00110110101001001000100100011100",
"01010101010011110111000000001101",
"01001010011001100111000101110001",
"01011100101001001111110000100000",
"01001110000100010101001000001111",
"01110101111010111000110010000010",
"01011010101011011010001101100110",
"00111000010100011100111100101000",
"00111011111001111100000110110100",
"01010110110110001011101111110111",
"01001011001001101000111100101010",
"00001010101100100010001111010001",
"00100101000101110000000011000101",
"00101100111110110001001001101111",
"00110110001100110100010010111111",
"01000111000100001011011101010111",
"01000011010000000111101000010011",
"00000001100011100101001111000111",
"00100000100001101111100101000000",
"01000100001000000101111111000111",
"01000001110010101001111101001100",
"01011010100110111010100110000100",
"01001101000011010010011110110011",
"01010011111010011000100100000100",
"01001001101011001110010011111101",
"00110011001011000111010010010101",
"00111001010100100001110110011001",
"01110000110001111000100101011111",
"01011000000111111101000010000100",
"01111101101111100001011001001101",
"01011110100110111111110000000100",
"01101010000010100011101100101101",
"01010100101111000001110101100011",
"01100111100000100100111111011001",
"01010011100000010010011010011001",
"00010000011111100001101001110101",
"00100111111111110000110011000110",
"00000000111000111101010101001010",
"00100000001010101100010101001110",
"01100111110011110101011000111111",
"01010011101000101110100010000111",
"01111011010100100011100111110000",
"01011101011001111111110010100111",
"00101001100101111101010100110010",
"00110100100010110110100001110100",
"00100010001010011111011010001111",
"00110000110100001001011110000011",
"00001011000111101011101101010101",
"00100101010010011001010100000010",
"00001000110000010100100000101001",
"00100100000111010100101000110000",
"01100011001100100100111011010010",
"01010001010101011010011010110001",
"01100001010100000100110100100000",
"01010000011001101110110000011101",
"00001001001111011000101100110010",
"00100100010111000100011110100001",
"01101001000101101110011000000000",
"01010100010001001000101110001111",
"00101000111000100110001110101101",
"00110100001010100011101010010000",
"00110111000100010000101100011111",
"00111011010000001011000111000010",
"00111110011001100101011000001101",
"00111110111100101101010001001001",
"00000101100001110101111111001101",
"00100010100000111010001010101111",
"00101100111111001001011110100010",
"00110110001100111100111101111100",
"01110110101110000010010100110110",
"01011011000110011000011011110111",
"01011100011000000001101111000100",
"01001101111011111000011000100110",
"00110111101011101011101101110011",
"00111011100101011000110100111110",
"00100011101100110011011110100101",
"00110001100101110111010101111110",
"00100011011100001101001100011011",
"00110001011110000100101111100000",
"00111001001111010000111100111010",
"00111100010110111111111110001100",
"01100111110100111001011101101100",
"01010011101001001001001000111111",
"01111110000011000111110010011111",
"01011110101111011010010010110110",
"00001101001001101001100000111111",
"00100110010011101000001110110111",
"00011011000000000000110000000001",
"00101101001101010000110101101111",
"01101110110101000000010111111110",
"01010111001001001011110100111001",
"00001010111001001010111010001100",
"00100101001010110001011010100110",
"00000101000010100100011100101111",
"00100010001111000010010110001101",
"01010110010101100101010111010111",
"01001010111010100011111000111101",
"00011011011000101100100100000001",
"00101101011100001111001101000000",
"00000101111011100001110001111001",
"00100010101011101001010010000101",
"00111110001001011010110000010111",
"00111110110011011111000100100011",
"00010110101101010000001011110001",
"00101011000110000011011100010111",
"00101111100001011111000110101011",
"00110111100000101111000000110011",
"01100000010011111010001010100110",
"01001111111001101000110110001011",
"00100001110100111011111001000110",
"00110000101001001010000101011011",
"00111000010001110011100111010101",
"00111011111000011101010111111010",
"01000011100000011111000101111001",
"01000001100000001111011111001011",
"00000011001001000000101101100110",
"00100001010011001110110110000011",
"01000001100001001100010100000111",
"01000000100000100101110011101101",
"00101100100110001101011101111001",
"00110110000010111101111011010100",
"00101100000001100110111100010011",
"00110101101110011000001101010011",
"01111000100101011101000000100111",
"01011100000010100111101001001011",
"01101010111111110010110110000110",
"01010101001101001011101001111000",
"00110001100011011100111011100000",
"00111000100001101011101000101110",
"00100101100100100110011111001001",
"00110010100010001110010011001010",
"01100001101101110101001010111100",
"01010000100110010010111100100000",
"00001101111011011110101010100100",
"00100110101011101000001000111111",
"01011101010000010010001100111100",
"01001110010111100101101110111100",
"00000101011010101000101001100001",
"00100010011101010000100100010011",
"00110001010111101011110110111111",
"00111000011011101100101011010001",
"00010110011111100011001001110110",
"00101010111111110001100011010010",
"01101101001111100010000111001101",
"01010110010111001001111100010011",
"00101111011010110011101001011111",
"00110111011101010110010011110001",
"00100011101001001100101010110101",
"00110001100100010011110001001001",
"00001000001111100010110111001111",
"00100011110111001010011000001010",
"00011110001111110100000001011101",
"00101110110111010100010100010110",
"00101110100010010111100101000001",
"00110111000001001010011011111100",
"00001101010010000111010011111110",
"00100110011000101000100001010100",
"01110100100101011001011000110101",
"01011010000010100101111110000001",
"01001001111011000100001001000010",
"01000100101011011110011001010110",
"00010011001101101001000101110111",
"00101001010110000011000001000001",
"00110010101110110100001001001100",
"00111001000110101101000111011000",
"01100000101000010100010100110011",
"01010000000011111010110011100001",
"01000010101111001000001100100010",
"01000001000110110101011001000001",
"00010011000010101110010011110010",
"00101001001111001001000011000100",
"00000010011101010000001101111010",
"00100000111110100111001001010000",
"01111011000000111011110011110111",
"01011101001101111010010011000010",
"01010110100011001101011001101011",
"01001011000001100100001111110100",
"00000101100110010000111011100000",
"00100010100010111111100000101011",
"00111100100010001000000111111111",
"00111110000001000010111101111001",
"00000011001001011010110111100100",
"00100001010011011111001001000010",
"00110001100111110111110111110100",
"00111000100011101110000110001000",
"00110101000111100101001000100110",
"00111010010010010101001000101101",
"01101110001001001101101101101011",
"01010110110011010110111101001000",
"01100011001011010100110011010100",
"01010001010100101010000100101100",
"01011010101100001011100111101111",
"01001101000101100110011100010101",
"01001111110111000010111000100111",
"01000111101001111110000011001110",
"01110001000110110011011101111001",
"01011000010001110101011001101011",
"00110111111100011101110100101011",
"00111011101011111111001101010100",
"01010101010001101011100010001001",
"01001010011000011000110010100110",
"00100010011110011111010100111000",
"00110000111111001111010111111101",
"01001110011100000000111110100001",
"01000110111101111110011100000110",
"01000010100001001101101001010110",
"01000001000000100110011101100100",
"01010001111001010010111110010111",
"01001000101010110100011011100110",
"01110010000101001101101001010111",
"01011000110000110011010101011101",
"01001010110000110000100000100101",
"01000101000111100000000000001110",
"01110000001001000110111111110101",
"01010111110011010010110001001000",
"00100000100111100101001110011000",
"00110000000011100101101110100101",
"01011000000010110111110100100011",
"01001011101111001111011111110111",
"01100100101110100000011000101010",
"01010010000110100100111011110010",
"01101010100010101001010111011011",
"01010101000001010011000000000100",
"01101011010000100000111010011010",
"01010101010111101110001100001111",
"00010111011101010100100001110110",
"00101011011110101001010110010000",
"01001011001010111101101100001110",
"01000101010100011011111111111110",
"00101101111111101001000110111101",
"00110110101101001000001101000101",
"00101010100000000010110101101000",
"00110101000000000001011010110001",
"01001101101000001101111010001000",
"01000110100011110111111100011111",
"00101001000000100100111010110100",
"00110100001101101010010011000101",
"00000001000011010000001111010100",
"00100000001111011111111111100001",
"01010011001110011110110101101001",
"01001001010110100010101100010101",
"01100101100010101101000010110011",
"01010010100001010100110001000111",
"00000100001100101011000110111000",
"00100001110101011110000111101010",
"00000100110110010110101101011101",
"00100010001001101101001010000001",
"00011010101010010010001011011001",
"00101101000100110010001100101101",
"01110010010101111000110100100011",
"01011000111010101110100000011010",
"01101000000001101011100000110001",
"01010011101110011011010111000000",
"01110101010110011101110011001000",
"01011010011011000010100110100001",
"01000010001100111011101101001011",
"01000000110101101000000010011110",
"01011001001000011110111110101010",
"01001100010010111001101101001011",
"00101101010010111011100111110011",
"00110110011001000101111101010100",
"00010111011110100111001111010100",
"00101011011111010011011000000101",
"01111011100110111110010011100011",
"01011101100011010100001010011011",
"01111011101110111100100110010101",
"01011101100110110000100110111011",
"01011001111111110100111000101010",
"01001100101101001100011000000111",
"01001101100000010001010001111010",
"01000110100000001000100111110010",
"01101101110100001010001111101100",
"01010110101000110110101101101001",
"00100100110000100101011001010000",
"00110010000111011011011111110110",
"00111101101001011000010001101111",
"00111110100100011000111000001011",
"00001110011011101111011110000100",
"00100110111101110101011000111011",
"01111100110011011101001101110011",
"01011110001000100101000001001011",
"00100010010111111000101010011001",
"00110000111011110011100010000110",
"01111000111110011000110101011111",
"01011100001100101011100110100011",
"01101000000011111110001000001110",
"01010011101111111110110000000111",
"00111001110101001101001100001111",
"00111100101001010000110011010001",
"01000100001001010110100001101110",
"01000001110011011100011100010001",
"00010110000011100111001111001011",
"00101010101111101111011100100101",
"01100100010101010000000001111000",
"01010001111010011000001101101000",
"00010001110001100100011011110110",
"00101000100111110100111100110011",
"00111111000100001100001001111111",
"00111111010000001000000101111101",
"01100101011000100000010001001100",
"01010010011100001000101010101011",
"01100101000000000011010001011111",
"01010010001101010010100111110110",
"00100100100110111001001100110011",
"00110010000011010001110110010100",
"01101001100101001011011000000100",
"01010100100010011111011110101000",
"01101001110110011001111110111100",
"01010100101001101110011010011000",
"00111111010001001011011000001100",
"00111111011000000110011111101110",
"01011011111011000100001100101000",
"01001101101011011110011010101011",
"01010001111000000101011111101110",
"01001000101010010111010100110101",
"00110100100111101001001011010101",
"00111010000011100111100000001111",
"00011110000111111111111001110011",
"00101110110010100110000111000111",
"00101011000000100100011110011000",
"00110101001101101001111111001010",
"01100001111010100100110011001000",
"01010000101011010010110101100101",
"00110101100110100111001001000111",
"00111010100011001001101001001111",
"00100110100111100010110001111011",
"00110011000011100100101000001110",
"01011101101001100001011001011101",
"01001110100100011100111000100111",
"00001111100110011100000001110001",
"00100111100011000100100101000100",
"01110100000111110100000011110110",
"01011001110010011110100111001010",
"01001011011101101011101001001001",
"01000101011110110101001000110010",
"00110100010111000001011011000001",
"00111001111011010101110111000100",
"00110001110001001100010101100101",
"00111000100111101011010000000010",
"01011001111001011011000111001110",
"01001100101010110111011110000111",
"00110001001010011110101000110101",
"00111000010100001000111111101110",
"01010100001001000100111111111111",
"01001001110011010001100001010111",
"01010010110111110011111100101101",
"01001001001010010000101100001100",
"00011001001110011100110001000011",
"00101100010110100001011110100010",
"00001101111110010010001100001110",
"00100110101100101001001110001110",
"00010111000001001010011110011011",
"00101011001110000100100000000100",
"00101111010010000100000000001110",
"00110111011000100110101001101000",
"01110010010011100010001110000110",
"01011000111001011011100001110100",
"00101000110010101110111010010010",
"00110100001000010010101100100010",
"01101110010110010000001010001101",
"01010110111010111011001100111011",
"01010111101100000010011111010010",
"01001011100101100010100011011100",
"00001101110010110010001011110001",
"00100110101000010011111111101100",
"00010010111101001001010111000000",
"00101001001100001110111111111111",
"01000001010001001101110111010111",
"01000000011000000111111010100000",
"01110111101001001100001010101110",
"01011011100100010011100011000000",
"01010010001110010100101111001101",
"01001000110110011100110000101111",
"00011101001100010010000011111111",
"00101110010101001111000110010001",
"01001001100001010001101010011100",
"01000100100000101000011011101011",
"00000110110101111101111010100010",
"00100011001001100011101000001000",
"00111011010100010001111101110010",
"00111101011001110110000010010101",
"01110100100001110110001000110100",
"01011010000000111010001111011010",
"01101000110000100010101101101010",
"01010100000111011010011010001100",
"01110000111010111001000110111001",
"01011000001011011010010101010010",
"00011011001001011000111010110000",
"00101101010011011101111011011100",
"01000110011010000100000111001000",
"01000010111100111101011011110011",
"00000000100001010101001000101010",
"00100000000000101010001000100101",
"00001111010001001100111110100110",
"00100111011000000111011010001000",
"00010001110111101111110000010001",
"00101000101010001111000110100001",
"00110100111000010110100011101100",
"00111010001010011101110000110000",
"01000001000010011001010100001011",
"01000000001110111010110000110101",
"01101011110001001010110111011111",
"01010101100111101010101010000110",
"01100110000010110101001100100001",
"01010010101111001101101110000000",
"00010101001011011110010100001010",
"00101010010100101111110110011000",
"00111110101000111110110100001101",
"00111111000100001101101001111100",
"01111111010001010001111101100100",
"01011111011000001010001111111100",
"00100011001001110000100000011001",
"00110001010011101100100011111110",
"01010101101010001001010010101000",
"01001010100100101110010101001000",
"00101110100011010101111101110010",
"00110111000001101000010100110101",
"00010101011101010010101110011111",
"00101010011110101000011011010100",
"01111110011100111000001100111010",
"01011110111110011010110110100001",
"00011100111001100110000111111111",
"00101110001010111011100100111110",
"01101101001001010101001101110010",
"01010110010011011011101000000011",
"00001100001111101010011000101100",
"00100101110111001110101111010010",
"00101111110110101111011111000000",
"00110111101001110110101001001111",
"00101110011010100011000101001001",
"00110110111101001101101010000101",
"00000011111000110110100011011010",
"00100001101010101001110010100110",
"00000010000101000100001110001101",
"00100000110000101101001001100100",
"01001011100110110101001001001000",
"01000101100011010000000000100000",
"01001101011010001000001101110110",
"01000110011100111111100101101011",
"00001000111011000010001000101111",
"00100100001011011101101010001000",
"00000110111011000111000110111010",
"00100011001011011111011111001110",
"01000001111011111110010110101010",
"01000000101011110011101111010000",
"01110001101011100100110110011001",
"01011000100101010101111000110100",
"01110111110110000000001101110011",
"01011011101001100100100000110100",
"01011101000101010111010001011010",
"01001110010000111001101000111111",
"00111000000101101000111101100001",
"00111011110001000101001100011110",
"01111000010111010101010110011101",
"01011011111011100000100101111000",
"01101100010110100100010000000000",
"01010101111011000110000110001100",
"01001001111101011000101101110011",
"01000100101100010100100011001000",
"00101101001111101011111010001001",
"00110110010111001111100111101111",
"00101101011000111101100100001100",
"00110110011100011000001110011001",
"00110101101110100011100101010010",
"00111010100110100110010000101001",
"00010011010010100001000110101010",
"00101001011000110111000100001010",
"01000010100100011011111000010110",
"01000001000010001001010101011110",
"01110100010111100010011001011111",
"01011001111011100111100110011111",
"00010010100011110011000100001110",
"00101001000001110110001000000101",
"01100101101110001100011000101111",
"01010010100110011100101000000010",
"01001010000001101011101100001000",
"01000100101110011011011110110110",
"01000001000111001001000010000000",
"01000000010010000011001101111101",
"01111011001011011111000111001111",
"01011101010100110000010101010111",
"01001000011110100011111001000010",
"01000011111111010001101011101111",
"01011110000000101111001010000000",
"01001110101101110001011101101100",
"01101000010100110100010101000001",
"01010011111010001000111111110111",
"01010100101110001110010001101110",
"01001010000110011101011010011000",
"00001101110111011110101001000000",
"00100110101010001000100111000111",
"00010110101111010111011010001010",
"00101011000110111011101001101010",
"01011000100111000100110101001000",
"01001100000011010111000111100000",
"00001111111100100010110111001101",
"00100111101100000001000010100110",
"01100010010110001100100011010010",
"01010000111010111001001111011110",
"00100110000001001101000010111110",
"00110010101110000110010010010100",
"00011000110111100100111111111100",
"00101100001010001011000001100100",
"01101001010001010011101010001100",
"01010100011000001011001101110101",
"01100111111101001011011001101001",
"01010011101100001111101111001110",
"00001010100011001001110110010101",
"00100101000001100010100011011001",
"01100001000111010011110111111111",
"01010000010010001010001001001101",
"01000101000010100010101011000011",
"01000010001111000001001000110110",
"01000010101000110010110011110111",
"01000001000100001000010110000100",
"01011001011110101001001110011100",
"01001100011111010100011000010101",
"00110001011001000110111011000100",
"00111000011100011101001011100101",
"00001100100110001011100001101010",
"00100110000010111101000010011101",
"00000110101110010101001000100110",
"00100011000110100000010000110111",
"01011110110010000100011111010000",
"01001111001000000001110010110110",
"01000010010100101111000110111100",
"01000000111010000110000111111010",
"00011010000000110110001111010000",
"00101100101101110110011010010011",
"00100001010110100000010111100110",
"00110000011011000011111111101000",
"00110110101100010001100000011100",
"00111011000101101000111100100100",
"00101100100100101001010011011111",
"00110110000010001111100111011101",
"00000111000100101100110000010110",
"00100011010000011101101100010111",
"00000000101101111101001100100100",
"00100000000110010110010010111100",
"01101101101011110010010101011111",
"01010110100101011011101010001011",
"00000010010000001011110111100101",
"00100000110111100010000101011110",
"01001001001100100001000101100110",
"01000100010101011000000111100011",
"01001011101100100001011111011111",
"01000101100101101111101110110100",
"01101010100101000000001100100110",
"01010101000010011010010010010110",
"00011101111010101111010111010101",
"00101110101011010110101111010011",
"01011001100100000000001000011111",
"01001100100001111100010010110101",
"00000001010100010111100110110000",
"00100000011001111001001001111100",
"01110110100001110100001100011101",
"01011011000000111001010010111011",
"01101001100000100010111111101100",
"01010100100000010001011011000101",
"01100011101010100100001010000010",
"01010001100100111010000000011001",
"00011100100011000001001111011100",
"00101110000001011110011100010110",
"00000010011000000111111111101000",
"00100000111011111011101110100100",
"01001100111011110111110100001110",
"01000110001011110001010110010111",
"00000100100000001100101001000101",
"00100010000000000110010011111010",
"00001100111011010001110101111110",
"00100110001011100011011011110010",
"00101110000011001011101100001101",
"00110110101111011100111011010101",
"01001001100010101111010100001000",
"01000100100001010101110110111000",
"01001111100100000100101001110101",
"01000111100001111110011011001010",
"00000111100001110100111010101001",
"00100011100000111001101001011001",
"01111010111011110110001111001100",
"01011101001011110000110001011011",
"01011100001010010000001011011111",
"01001101110100000000000111000011",
"00001110010000001010000011001111",
"00100110110111100001000010011011",
"01011001101101111010101110011100",
"01001100100110010101010000111101",
"00011110011110111111010010011011",
"00101110111111011111100000111101",
"00101000010001000000010010100000",
"00110011111000000000001010100100",
"01111011000100011011000110000011",
"01011101010000010010000000101001",
"01010101001011010000110010110111",
"01001010010100100111101000110011",
"01010100110101101001100101111111",
"01001010001001011011110010101010",
"00000010001001000111110110011001",
"00100000110011010011010011001010",
"01010101111001001101111111011011",
"01001010101010110010100100011000",
"01000010100001011011111011011110",
"01000001000000101101011101011100",
"00000100011001010011101101111110",
"00100001111100100011111100101010",
"00011111000101101111000101000010",
"00101111010001001001001011100100",
"00001110001101111101011010111110",
"00100110110110001111000010000010",
"01101110111110010011111010100100",
"01010111001100101001110101110001",
"00111101000000011110011100010111",
"00111110001101100101110000011001",
"01100111110001111101100011011101",
"01010011100111111111000001010111",
"01110000010010101011100001010100",
"01010111111000111100111011000010",
"00110011100010010010101000110100",
"00111001100001001000000011010010",
"01010001010010100000100011001010",
"01001000011000110110110000001011",
"01010011111101001111101011010110",
"01001001101100010001010010001011",
"01010000000101010011111000010000",
"01000111110000110111011010110110",
"01010011101010101000100010110010",
"01001001100100111011111010000011",
"00100000111001000111011111100100",
"00110000001010110000001000110011",
"01010100100101100000100001010101",
"01001010000010101001010000111111",
"01100000100101111010011000110000",
"01010000000010110101001011011101",
"01001110111100010011001011110001",
"01000111001011111011010101011110",
"00011110001000001111110101011110",
"00101110110010110000001011000000",
"00110000001001111111000010100101",
"00110111110011110101100010111111",
"01010110011110001000000110011010",
"01001010111111000011100110101100",
"00011001000100000110000100101010",
"00101100010000000100000010111011",
"00001100010100001111001110000100",
"00100101111001110100100001000101",
"01100100101110010010001001101010",
"01010010000110011111000001011111",
"01110010110010000000110011000111",
"01011001001000000000010100011100",
"00101010110011001110100000100000",
"00110101001000011111001101100111",
"00001100111111010010011100001010",
"00100110001101000000001010000000",
"01101101110110011011111001001010",
"01010110101001101111001001001111",
"01100001110100111100000010001001",
"01010000101001001010001000111100",
"01101111111111100011101111100011",
"01010111101101000110010011010010",
"01010101110111101101010010110011",
"01001010101010001110001010110111",
"00100100010110010111111101100111",
"00110001111010111111011011111111",
"01110100011000110111011101100001",
"01011001111100010100111111010001",
"01110100111101011100010111110101",
"01011010001100010101110111100101",
"00110010100100010101011000100101",
"00111001000010000110010010100000",
"01100011010111001011011000000101",
"01010001011011011011001110010111",
"00110001111101111010110100001100",
"00111000101100100000110101010001",
"00011010010110010010111100000011",
"00101100111010111100101101011111",
"01010011101001110110111001011001",
"01001001100100100110010011010101",
"01100101100000001101011101000000",
"01010010100000000110101101110011",
"01101011101000110011011111001101",
"01010101100100001000101001010001",
"00100111100111000110100100101111",
"00110011100011010111111001111111",
"00110101100101100001010101010001",
"00111010100010101001101000111110",
"00111111010011011100000001111111",
"00111111011001011000000101000000",
"01001000100000001110000100010011",
"01000100000000000111000001010111",
"00001010001011000001110110100110",
"00100100110100011110100010011110",
"00011111111001010110011010110000",
"00101111101010110101101101111011",
"00010111011100100001010000000100",
"00101011011110001111000100011000",
"00101000010011010001101100000100",
"00110011111001010010010011100010",
"01010000000011010101011101010101",
"01000111101111100011100000011011",
"01101101111010101001010110011110",
"01010110101011010100100001001110",
"01000001010111010111110000101111",
"01000000011011100001111000110100",
"01011100010111100100101011011010",
"01001101111011101000110100110011",
"01010010101000111011100000001000",
"01001001000100001100001100001101",
"00110100001001011000100011110110",
"00111001110011011101101101001101",
"00000111001010110011001011111010",
"00100011010100010101100101010011",
"01011111101000001101111100010010",
"01001111100011110111111101011100",
"00100001111111110100011101000000",
"00110000101101001100001110010101",
"00000111001001010010011111010001",
"00100011010011011001111011011100",
"01000001011101001001111110011011",
"01000000011110100011111101000000",
"00010001111111011000001100100011",
"00101000101101000010001100111100",
"01011101000000111111110010000100",
"01001110001101111101000100000111",
"01100101110011100001111100000011",
"01010010101000100110111000010100",
"00000110011000001111101010000100",
"00100010111011111111110100010011",
"01010001111110011100001001111001",
"01001000101100101100110010100111",
"00011000010111110111010100101000",
"00101011111011110010110100001101",
"01101001101111011011000010001001",
"01010100100110111101001000111110",
"00000011111100010110111110000101",
"00100001101011111100101101101110",
"00110010101110001010010000101011",
"00111001000110011011101111011010",
"00111101011001010001111011100010",
"00111110011100100011000000001100",
"01101001011100100100011011000110",
"01010100011110010000101100110001",
"00011110010110111101101111111000",
"00101110111011010011111000001111",
"01100101000000011000100000010001",
"01010010001101100001100101011011",
"00011111000010000101110000010111",
"00101111001110101101011001001001",
"01011101101010011001110001111000",
"01001110100100110101100000001100",
"00101101100000100110100100100100",
"00110110100000010011001100100001",
"00101001001101000111100110111101",
"00110100010101101111001000100101",
"01111101100011110000001100101000",
"01011110100001110100110001010000",
"01000100111101000111110100101000",
"01000010001100001110011100011001",
"01010001100000011001010011000010",
"01001000100000001100100111000010",
"01001101100111000101101001111101",
"01000110100011010111011111011010",
"00110010110111110001001011000110",
"00111001001010001111101000111011",
"00010010110111110001000011110001",
"00101001001010001111100110001001",
"00101001111110101010010101010111",
"00110100101100110001110111001001",
"00000101100000101100101011001111",
"00100010100000010110001101111001",
"01000111000001001001100111100111",
"01000011001110000011111001111111",
"00110001001001011101100001010001",
"00111000010011100000110010011111",
"01100101001000111010100111100001",
"01010010010011001011000010010000",
"01101001000000111110000100100111",
"01010100001101111011110111111000",
"00111000010010110000000000100011",
"00111011111000111111011100010111",
"00100110100110000100100101111101",
"00110011000010111001110111001101",
"01111011000000010110010001001010",
"01011101001101100000000000110100",
"00010101010011101111110010100111",
"00101010011001100011000101010000",
"00001100011001100110100010000000",
"00100101111100101101111000000011",
"00000001011000100101111011001110",
"00100000011100001011101011001111",
"01100111010010001011111100100001",
"01010011011000101011001000110100",
"00100100110001011101110110101000",
"00110010000111110010010011011111",
"01101011001000000000111101010111",
"01010101010010100110110001110101",
"01101011001110100010111010100110",
"01010101010110100101000101011000",
"01010111011111101000000111010100",
"01001011011111110100000010100010",
"00101000100001010010111000111001",
"00110100000000101001000010001000",
"01010100101011000111010101101100",
"01001010000101001001001101011010",
"01110101110110100101110111001100",
"01011010101001110010111101101010",
"00001101100001101011011001001010",
"00100110100000110101000000101010",
"01110011101101001101000110000011",
"01011001100110000010001001001101",
"01010011100000111111101001000100",
"01001001100000011111100100111100",
"00111011000010010001111101101110",
"00111101001110110101101111101101",
"00011100111010010100101101000001",
"00101110001011001100111000011110",
"01010001000100101111110101101100",
"01001000010000011111101110101001",
"01101110011010101110000000000011",
"01010110111101010011010111001011",
"00011110101011110101011111101010",
"00101111000101011101000000100101",
"00110010110111001010111101011100",
"00111001001010000001001000001001",
"00000001010010011111000011110100",
"00100000011000110101111010100000",
"01001000101010011111110101000001",
"01000100000100111000001000001111",
"00111000010111110111101000101011",
"00111011111011110010111110111011",
"01001000010011101000101011011011",
"01000011111001011111001000000000",
"01111001110011111101010110010011",
"01011100101000110001101010000101",
"00011101100000110010010000001101",
"00101110100000011000111110010110",
"00110001010100100110110000000010",
"00111000011010000001100001000110",
"00110010000110101101010110110110",
"00111000110001110001011110011011",
"01000100000110110110110110001010",
"01000001110001110111100100011111",
"00101100010100111101000001001100",
"00110101111010001101110001110001",
"01000111011010011101001001011101",
"01000011011101001010100011100000",
"01010000100000011101011000001010",
"01001000000000001110101000101110",
"00101101101101100010111100011010",
"00110110100110001011010100011000",
"00101110101100101001000101111110",
"00110111000101110010111100111001",
"01110101010001111011001110110010",
"01011010011000100001101100000001",
"00011000110101100011111001110001",
"00101100001001011001100101111110",
"00011001111011001100000000100101",
"00101100101011100001010010100100",
"01001100110001100011010110000110",
"01000110000111110100100000110010",
"01000001010110110110110010101010",
"01000000011011010000000111111001",
"01101110100110010011010110010001",
"01010111000011000000100111011011",
"01000010101000001001001101010011",
"01000001000011110101110110001111",
"01001110111000100010001011110100",
"01000111001010100010001000111010",
"01100010010011100000011100010101",
"01010000111001011010100010011011",
"00010110001001001000110110010111",
"00101010110011010011111011000100",
"00001001111010110100001001100010",
"00100100101011011000100000010001",
"01111111001101110101001001010110",
"01011111010110001010001001010100",
"01100111001101111000101100000100",
"01010011010110001100001111001110",
"00001001111010001101111011111000",
"00100100101011001010011000000000",
"01101101101000100011001001011001",
"01010110100100000001011001011110",
"00000101111001101110001011101110",
"00100010101010111110100101000100",
"00111100110001011000111001010100",
"00111110000111110000010011110110",
"01101110111011000010001101001101",
"01010111001011011101101011110001",
"01001110100100001110000000101111",
"01000111000010000010110100111011",
"01110101001001010000100010000000",
"01011010010011011000101101011100",
"00110111001110101010111000101000",
"00111011010110101001110000001101",
"01001000011000001011010111000010",
"01000011111011111101100001100011",
"00010010101010000010110010001101",
"00101001000100101011011111100101",
"01101000100011010001101000101010",
"01010100000001100110010000111010",
"01111010011110111000101101111000",
"01011100111111011100001100111010",
"01010110110000111001101000010111",
"01001011000111100011101100100001",
"00010100111000001110101001110110",
"00101010001010011010110010000100",
"01000001111001010101110111010110",
"01000000101010110101100000101101",
"00100111010001010111000000100001",
"00110011011000001101000111111000",
"01000010100101110001100110010000",
"01000001000010110001001000110110",
"01110000100101111110111101010100",
"01011000000010110111010001110011",
"00011100100011010010001111010011",
"00101110000001100110100011010100",
"01011011011011010101100000000001",
"01001101011101100111111011010101",
"00001010100001001010111101111001",
"00100101000000100101001001011000",
"01101001010100110101100101011010",
"01010100011010001001101100000110",
"00011100110010001100010010101011",
"00101110001000000100111010010110",
"01111001000111011110010100001011",
"01011100010010010000110011000010",
"00101011111100111110110010101101",
"00110101101100001011001011001100",
"01101011101010101110011110011111",
"01010101100100111110011110011100",
"01011011011010111110110000100000",
"01001101011101011100000110010111",
"01000010000110000111101001000100",
"01000000110001011001001000100111",
"01110101100101100010101000000001",
"01011010100010101010001111001011",
"01011010101000110011111001110110",
"01001101000100001000110101000100",
"00101001010100000000010101001000",
"00110100011001101100010001000111",
"01111111011111110000100011111001",
"01011111011111111000010001011110",
"01001000010001010111000011001111",
"01000011111000001101001001011011",
"00101111001101101110100000110110",
"00110111010110000110001110010111",
"00111100010001001001011101001101",
"00111101111000000101011001100011",
"00110111001100011001010000011100",
"00111011010101010011011010111001",
"01111101110001111100100001100110",
"01011110100111111110100111000000",
"00110001011010011001111111001101",
"00111000011101001000111001101011",
"01101110011011000100001001000100",
"01010110111101011110111001110001",
"01000110001010000111111000101000",
"01000010110011111011000000001000",
"01000100000100011100110001011010",
"01000001110000010011000111110011",
"01010110111110010101110001101110",
"01001011001100101010100000011100",
"01000000101001000000100110100001",
"01000000000100001110011100011011",
"00011010110101010110011001110001",
"00101101001001010100010111101110",
"01101011110110100100011011100100",
"01010101101001110010011010100101",
"00000010100010010110011101110111",
"00100001000001001001111001100110",
"01000010000110101101011010010010",
"01000000110001110001100000101001",
"00101110011100010110000001110100",
"00110110111110001001010010110011",
"01110011001000010101011011001011",
"01011001010010110011101100011011",
"01011110101001111111101001100110",
"01001111000100101010001000000100",
"00001001110111101011100001110101",
"00100100101010001101100000000010",
"01111101101001100000011001000101",
"01011110100100011100011100010110",
"01000111111110110101001111000000",
"01000011101100110101110000010000",
"00100110101001110111110100100000",
"00110011000100100110101101001011",
"01110110110000111110101101010000",
"01011011000111100101101111111000",
"01110011111011110100000001101101",
"01011001101011101111111101101011",
"00010010010100100110010010111111",
"00101000111010000001010001000100",
"01010010001011111101011101110000",
"01001000110101000010101100011101",
"00110110000001111011101010110001",
"00111010101110100110011110010111",
"00000111111010001000111011000000",
"00100011101011001000100001000000",
"00101100110100110001010111100110",
"00110110001001000101111111011001",
"01011111010101111011111111111010",
"01001111011010110000001111001100",
"00000111011001111001011110111001",
"00100011011100110111110110011110",
"01110101000110001000011010110101",
"01011010010001011001101000110101",
"00001110100011101010100000110000",
"00100111000001110010000101000001",
"01000011101011000010111100000110",
"01000001100101000111010100000100",
"00101100010010100001101011010001",
"00110101111000110111011000110001",
"00001100010101100111000010010110",
"00100101111010100100110011011001",
"01110101000101011100111011010100",
"01011010010000111101010101101011",
"00011010101101100101110100010101",
"00101101000110001100100001011100",
"01010010011111101110111010111111",
"01001000111111110111011100111010",
"00111001001001111001101100101110",
"00111100010011110010001111110101",
"01110001101011111011100110000011",
"01011000100101011111100111010001",
"00010011001000101111100001100000",
"00101001010011000100000101110011",
"01010011111111010000000110100000",
"01001001101100111111010100110010",
"01011101100010100000000001100111",
"01001110100001001110100000011111",
"00010101101011000101111111010111",
"00101010100101001000101000001110",
"00010110000101111101100000110010",
"00101010110001010010100100001011",
"00001011111110110110000011011011",
"00100101101100110110000010111100",
"00001000110011011011011010100010",
"00100100001000100100010011101110",
"01110100101111111101001010011000",
"01011010000111001011000111100101",
"00010101110110100001100101010000",
"00101010101001110001010100110001",
"00000110011100111011110011100111",
"00100010111110011100101100110000",
"00111100101110110010011001011000",
"00111110000110101100011001001010",
"00111100100000011001011001110000",
"00111110000000001100101010011000",
"01111101001101111010100000110111",
"01011110010110001101010100001100",
"00110000101010100110011011000101",
"00111000000100111010111111001111",
"01001110110100111111101100101111",
"01000111001001001011100100000111",
"01001111011001110111111110100111",
"01000111011100110111000011110110",
"01100110101100100010000101110111",
"01010011000101101111111111000101",
"01010110101111001000100111101111",
"01001011000110110101100100001110",
"01111100001110101001010110001101",
"01011101110110101000110110100100",
"01000110000010011110000101110001",
"01000010101110111110000001001010",
"01011110001001000010000110101000",
"01001110110011001111101101101001",
"01110001010100110001110001000010",
"01011000011010000111100101100101",
"01010100100110001000100110100001",
"01001010000010111011101100110001",
"00100001110100000101000010101110",
"00110000101000110100101011001100",
"00011101100111010011011100010011",
"00101110100011011101101110000001",
"01100000111011101111101000111000",
"01010000001011101110010110111101",
"00010110111001100001111110000010",
"00101011001010111010000001110101",
"00111000010100111001010000101000",
"00111011111010001011101101100000",
"00110011011011011110100011110111",
"00111001011101101100101000001111",
"01010000000011011011101010110001",
"01000111101111100111101011101011",
"00101010000000110100110110101011",
"00110100101101110101011100011101",
"01000110100100001110000101010111",
"01000011000010000010110111000110",
"00100100000010101011110001010001",
"00110001101111000111010100101110",
"00000111100011010100111000010010",
"00100011100001100111110011110000",
"01011100001111010100000100101110",
"01001101110111000001110010011010",
"00111010001000101001010010000011",
"00111100110011000000001011010101",
"00010011100010001010111011101101",
"00101001100001000100010100111001",
"01100101000010101111011111010000",
"01010010001111001001110110010010",
"00101110111000100110011100011100",
"00110111001010100011101111011011",
"00101001011000101100100000111101",
"00110100011100001111001011011000",
"01101011011111101011010010111000",
"01010101011111110101101000100101",
"01101011100111011000110101110100",
"01010101100011100000001001110101",
"01100101111001000101111010101101",
"01010010101010101111100011000011",
"01101000101101100101110011101111",
"01010100000110001100100001001100",
"00011100010001111111010000111010",
"00101101111000100011111110000110",
"00110100101110000101100111011100",
"00111010000110011001110011101000",
"00111000000111011101110010010111",
"00111011110010010000011101100000",
"00000010111110100001010110110001",
"00100001001100101110101001101110",
"00001011011101001110001111001011",
"00100101011110100110001000011111",
"00110100010110000111001000100100",
"00111001111010110110010011000001",
"01001001000000111111011100100010",
"01000100001101111100110101000111",
"01101001100110010000010101110011",
"01010100100010111111001111011011",
"00100101101010111000111001100111",
"00110010100101000010111110110101",
"00011101100111001000000011000011",
"00101110100011011000100100101001",
"00001011011010010101011000100010",
"00100101011101000110011111011001",
"01000011010010001100010101111010",
"01000001011000101011010111001001",
"01111110100010110111101011111011",
"01011111000001011001110111110000",
"00100010010011110111010110100100",
"00110000111001100111010010001100",
"01111011100111000101100110100011",
"01011101100011010111011101110111",
"00110001111110010110001111110010",
"00111000101100101010101011001101",
"01110010010111010011000001010101",
"01011000111011011111010101101011",
"00100101100111111010011101001110",
"00110010100011101111010000001100",
"01111000100010100100010101001001",
"01011100000001010000100101000110",
"00010110011001111110110010100110",
"00101010111100111010101000111110",
"00101101001011001111010101100001",
"00110110010100100110110000000001",
"01010100110001111000011001110111",
"01001010000111111100111101011010",
"01010000100010101000000100101010",
"01001000000001010010011000010010",
"01000000101101011010010001001110",
"01000000000110000111101011100001",
"00111001110100100111111001001000",
"00111100101001000010010011000110",
"01111111011011001110100001000110",
"01011111011101100100010011001001",
"01101010000110000110110010001100",
"01010100110001011000100101000011",
"00100101010100010011001100000000",
"00110010011001110110101101100110",
"01101011000010100111010110111010",
"01010101001111000100010100110110",
"01001111111111001100101100111001",
"01000111101100111110000111011000",
"00001110000001111000111111101111",
"00100110101110100100101000110111",
"00000111010100100110100111110100",
"00100011011010000001011100100100",
"00000100101101010010010100010110",
"00100010000110000100010101110010",
"01000110001001010110110010000110",
"01000010110011011100100110011110",
"00001010010011000111111110100101",
"00100100111001001100111000001000",
"00010000001010100000100011100001",
"00100111110100001010001011000000",
"01111010011111011101111010101011",
"01011100111111101110111011000011",
"01010011010100000111011011000111",
"01001001011001110000001100110011",
"01111001110000110000111001010101",
"01011100100111100000001010010000",
"00100000001010010110110100010010",
"00101111110100000100001100010011",
"01110000111011001111011110001011",
"01011000001011100010100100000001",
"00000101001011000110010001110111",
"00100010010100100001001111001000",
"01100011011100100011001010001100",
"01010001011110010000000011001010",
"01101111011110000111001010000110",
"01010111011111000011001000000101",
"00100111011110111101101000011011",
"00110011011111011110101011100010",
"01011111000011101000110000101111",
"01001111001111110000011101111110",
"00100001011100011101011001111001",
"00110000011110001101000101110001",
"00011001110110010000101001110001",
"00101100101001101010110101001111",
"00000100101011100011001101111110",
"00100010000101010101001100000100",
"00011001111111000001101111000010",
"00101100101100111010001101011111",
"00110000010000001111011100010111",
"00110111110111100100001001010001",
"00110001110110110010100011011111",
"00111000101001110111110100010101",
"01101110110000111010001000111010",
"01010111000111100011111001101100",
"00000000110010110111100001000001",
"00100000001000010110000111000101",
"01110010100100001100110100101101",
"01011001000010000010010001001100",
"00101000100101100010000010000010",
"00110100000010101001111101101000",
"01011100101010010011100110111001",
"01001110000100110010110100100000",
"01001101111001110101001110000010",
"01000110101011000001001100101000",
"01101011010000101101011001000010",
"01010101010111110101010110011011",
"00101100101001100000010011110011",
"00110110000100011100011010000010",
"01011011111011101110001101110001",
"01001101101011101101110101100111",
"01110010100101010100000000110110",
"01011001000010100011011110110011",
"00110001010110110010101000001001",
"00111000011011001101110111111011",
"00100010000101000100111111111000",
"00110000110000101101101010001100",
"01111100111000011011111111011100",
"01011110001010011111110011101111",
"01000001100001010011001011101010",
"01000000100000101001001011010101",
"00011100100100100010111010100011",
"00101110000010001100101000010000",
"01010000001100100011011010100011",
"01000111110101011001100000110101",
"00111011010010000100000100111111",
"00111101011000100110101100010101",
"00111100101110111001101110110101",
"00111110000110101111011011001010",
"01000001000111110010111000101110",
"01000000010010011101110111100001",
"01000000011101001010010110110110",
"00111111111110100100001001100000",
"00100000001011011100111001000001",
"00101111110100101110111111000101",
"00110000100101111010000010110101",
"00111000000010110101000001011001",
"01100111111100000111111111010010",
"01010011101011110111010000010100",
"01111111001111000101101001110001",
"01011111010110111001011001000100",
"01010010000010010111011100101110",
"01001000101110111001011111010110",
"00000001110010011000101001000011",
"00100000101000001001110101100110",
"00000011111010101000110111101111",
"00100001101011010100010101110111",
"01101100000001011001001011110000",
"01010101101110001110101100110010",
"00110010000010101000000101011010",
"00111000101111000100110100011100",
"00110101110001011011011011001110",
"00111010100111110001010100111111",
"01011010110010010011010100101010",
"01001101001000000111101101111010",
"00110010110101011111100110011100",
"00111001001001010111111011100001",
"00101000010101101000001111111011",
"00110011111010100101011101110010",
"00000011010111110101010110101100",
"00100001011011110001110000110011",
"00110011000011100101101000100011",
"00111001001111101110010111110010",
"00000100111111111011110110110101",
"00100010001101001110110110000001",
"01010001010001101010100100101110",
"01001000011000011000001111101110",
"00011110010100010011000001100101",
"00101110111001110110100111110101",
"00110001101001011100001010101000",
"00111000100100011010100101100011",
"00101101001101011000110010100000",
"00110110010101111001010110011010",
"00010000111001100111000010011100",
"00101000001010111011111010110000",
"01100011000000001110110010110001",
"01010001001101011010110000000010",
"01001111010010011101110010011000",
"01000111011000110101001100101001",
"00001101110010000011000001111000",
"00100110101000000001001101100001",
"00100100100001100001111110011011",
"00110010000000110000011010100101",
"01101011110111000000101100111011",
"01010101101001111101001101111110",
"01011101111110100110011100011011",
"01001110101100110000011110001011",
"01011111110011100110000011011011",
"01001111101000101000100000000100",
"00101000100101111010011011110000",
"00110100000010110101001100110101",
"00011111000110011001010101001010",
"00101111010001100100100100101110",
"00100000010000110000011010010001",
"00101111110111110111000101001001",
"01001000110001010111010100110001",
"01000100000111101111101011011000",
"01001111101100010011010111111111",
"01000111100101101001101111010111",
"00001000001100111000011001100011",
"00100011110101100110000100001010",
"01001000000000011100111110100010",
"01000011101101100100101110100010",
"00100001101110101010110100101101",
"00110000100110101001010000101000",
"00001001111111010001000010100110",
"00100100101100111111101010001010",
"01001011111011000101110110010001",
"01000101101011011111000001100011",
"00001101110000000100000000011101",
"00100110100111001101111010011010",
"00111100000001111001001000000001",
"00111101101110100100101110100100",
"00000001101100100001010001011111",
"00100000100101101111101000111000",
"01101000100010010111010101001000",
"01010100000001001010010100010001",
"01101110110111011000101110011101",
"01010111001010000110010111010011",
"00101010000010001001100001011011",
"00110100101110101111111110001110",
"01101011111010001100101011110100",
"01010101101011001001111010010100",
"00100001111010111110010111000000",
"00110000101011011100010001001000",
"00101111000010000101011000010000",
"00110111001110101101001000101000",
"00111101001011110111010000100011",
"00111110010100111110111100101100",
"01000000001111010001011000100110",
"00111111110111000000001110010011",
"01100000101011100001100010111000",
"01010000000101010100011110001011",
"01101010011001010000000011000011",
"01010100111100100010000000100000",
"01010001001000111000011011000010",
"01001000010011001001101010011001",
"01000011101011110000010101101001",
"01000001100101011010110011100010",
"00111001101011101101110101011011",
"00111100100101011001101111000000",
"01011110111010111011011100111010",
"01001111001011011011001100100011",
"01101000001101010010010100000100",
"01010011110101110101100000001100",
"00100101100010101110100010010110",
"00110010100001010101011110111110",
"00111100111001100001111001010101",
"00111110001010111010000000000101",
"01001000000000111000010111011111",
"01000011101101110111111001010111",
"01001110001000101000111110000110",
"01000110110010111111111110110011",
"01011011111111111011001110011111",
"01001101101101001110100111101111",
"01101000010001101000110001110001",
"01010011111000010111001110011110",
"00010110111010000000010010110111",
"00101011001011000101010100000101",
"00101011101100001110100110011110",
"00110101100101100111101101011110",
"01110000011110100001001011010100",
"01010111111111010000010011111000",
"01011110111010011101010001011010",
"01001111001011010000000011011110",
"01001101011010111001011011001011",
"01000110011101011001010100100001",
"01111010011101110010001101111011",
"01011100111110111000011111000000",
"00101010110101100011000111101011",
"00110101001001011001010010100110",
"01011011001010111101011011101001",
"01001101010100011011110101110110",
"00110110011111101011010101111100",
"00111010111111110101101010001000",
"00101100100010000100011001001011",
"00110110000001000001001010001111",
"01000011101101010100110000110001",
"01000001100110000101010111100001",
"00100101010111000100000100011001",
"00110010011011010111010010011001",
"01010110100100001101111010100110",
"01001011000010000010110010000011",
"00101111100111100001011100100101",
"00110111100011100100000001110101",
"01000111010010000010011011011001",
"01000011011000100101110000100111",
"00000101100110010011010010110110",
"00100010100011000000100101110111",
"01101100110011011000101101001000",
"01010110001000100011001111010100",
"00000111100001010011110011111111",
"00100011100000101001011111000110",
"01100110010001110100110101101110",
"01010010111000011110000100010101",
"01010111001100101000110000001011",
"01001011010101011100101101011100",
"01011000101010001100001111000001",
"01001100000100101111100111001011",
"00101001111101100101001011010111",
"00110100101100011001000010110100",
"00010000111000010110100101100110",
"00101000001010011101110001011110",
"00110111100101000111101011111011",
"00111011100010011101110001000011",
"00010010001010110111011111011011",
"00101000110100011000001101101100",
"00110110011011000101000111111100",
"00111010111101011111011010011111",
"01110100011110101001100101010001",
"01011001111111010100100011111000",
"01011010001011101111110110111011",
"01001100110100111010011110011100",
"00000100100011101110000110000010",
"00100010000001110011110001100100",
"01010000011110100100110011110000",
"01000111111111010010001001011100",
"01000010011101011000101000101100",
"01000000111110101011011100011110",
"00011011011101101110011000111010",
"00101101011110110110100010010010",
"01111100001010110011011010001111",
"01011101110100010101101110000011",
"00110010111011111001110100000000",
"00111001001011110010000101000100",
"01111010011000001011101010010100",
"01011100111011111101101011110110",
"01001001100101101100110101011010",
"01000100100010101110111100011110",
"00101101011001101100000001111011",
"00110110011100110000110001011101",
"00100101001101101110110001111111",
"00110010010110000110011000011111",
"00100100110000101010010001000011",
"00110010000111011101011110010100",
"01100011111001010111010111110111",
"01010001101010110110000100101111",
"01010001101111110011001011001010",
"01001000100111000111000010010011",
"01101000011101111111000001110100",
"01010011111110111110111111111000",
"00001001010000011011011100010000",
"00100100010111101011000011000100",
"00101000010100000001000101110000",
"00110011111001101100101100000110",
"00011000000101100000011110011010",
"00101011110000111111101010000011",
"01010000100010011101110111101010",
"01001000000001001101011110000011",
"00101101111010010100011000100110",
"00110110101011001100110000111010",
"00000100111000111001001011100010",
"00100010001010101010110001101001",
"01011000000011110001101011101001",
"01001011101111110110011100001001",
"00010100001100001001001110010100",
"00101001110101001001110001111111",
"01011100000101100001111011101110",
"01001101110001000000100110111111",
"00110000101101111101111010101011",
"00111000000110010110100110001100",
"00111110001001101110011001101011",
"00111110110011101011010000100101",
"01101100111101111000100001010100",
"01010110001100100000000000011101",
"01101000010011000101100110100110",
"01010011111001001011100011000101",
"01010000010100100101111001000111",
"01000111111010000001000010110011",
"00100011011000111101101001010001",
"00110001011100011000010001000101",
"01011100110001101111001011110111",
"01001110000111111001010000111110",
"00101010100000010101110000000010",
"00110101000000001010110110001011",
"00100111111100101011101111010011",
"00110011101100000100010000111111",
"00101101010000010011111111101000",
"00110110010111100110110000111100",
"01101100111101101110011000101110",
"01010110001100011100010111000111",
"01000011011010011010001000001101",
"01000001011101001000111110011000",
"00101001011011000111011001110111",
"00110100011101100000100110011010",
"00011111111001101000001100101110",
"00101111101010111100010110011011",
"00111101110010100101110010100001",
"00111110101000001111000100100100",
"01110011000000110100001111010001",
"01011001001101110101000000111100",
"01001101010011010100001110101010",
"01000110011001010011101110010110",
"01100011000000010100100100100001",
"01010001001101011110110100011001",
"00010111110001011110100000010101",
"00101011100111110010100100010000",
"00110001001100101011100110100001",
"00111000010101011110011010100110",
"00110100110000000111101111101011",
"00111010000111001111011011111111",
"00111010011101000111000010110010",
"00111100111110100010011101000001",
"01011101000100001000110101011100",
"01001110010000000101111000100101",
"00011000010100111110000000100011",
"00101011111010001110010100100110",
"00001010111111100100111010011100",
"00100101001101000110101101110111",
"00001010111110011101001110000010",
"00100101001100101101001011000000",
"00011101001101110111001100000110",
"00101110010110001011010110100011",
"01100011000011010110100110000101",
"01010001001111100100010001010111",
"00011111001010100110011100010111",
"00101111010100001101110010000101",
"01111001010011011001000111110100",
"01011100011001010110011101001001",
"00010011110001010100100000110000",
"00101001100111101110100010111001",
"01011101010100010100110110000010",
"01001110011001110111101000001111",
"01100110010001010001101001001000",
"01010010111000001010000100010011",
"01111100000100011010000111010111",
"01011101110000010001010111000110",
"00101101101000111010101111001001",
"00110110100100001011110110100010",
"00001001101010001111010010011001",
"00100100100100110000111100001111",
"01011000110110001001010011001110",
"01001100001001101000000000011101",
"01011000001001010000011111001011",
"01001011110011011000101011101011",
"00110001100110111011000001101101",
"00111000100011010010101011010101",
"00000110000110011101010010110110",
"00100010110001100111001000011011",
"01000101000110111110110111111001",
"01000010010001111100101101111001",
"01110101000001010101001001111010",
"01011010001110001011111010001101",
"00101111100001100100101100101101",
"00110111100000110001101111101011",
"01100101000000100111000100101000",
"01010010001101101011110011101001",
"00110010110011111010111100011100",
"00111001001000110000101101101101",
"00100010100010011000111011111111",
"00110001000001001011000101111000",
"00110010010011111011010011010010",
"00111000111001101001011110100001",
"00010101110100001111100000111101",
"00101010101000111000110001101011",
"00111010010011110111011100010100",
"00111100111001100111010101011001",
"01100011100000100110111001110011",
"01010001100000010011010111000010",
"01001010100100010111010000101000",
"01000101000010000111001010110100",
"00111010100011010100111110011101",
"00111101000001100111110110101100",
"00011101111101101101111100100101",
"00101110101100011100001100111111",
"00100111101000100000000110000100",
"00110011100100000000000010101100",
"01010010111000010010111111000001",
"01001001001010011100011010100101",
"00101000111101010010110111000001",
"00110100001100010010011011110001",
"00110010100110111101010100000111",
"00111001000011010011101101101100",
"01110000000110001010001011000111",
"01010111110001011010110001100100",
"00001100000000101001011101000111",
"00100101101101101101011110011011",
"01010001110001100011110000011110",
"01001000100111110100101011011000",
"01101001011001100011010010111011",
"01010100011100101100001010111001",
"00011111110001111101111101110111",
"00101111100111111111001011111011",
"00101111000101111000100110100000",
"00110111010001001111011000000010",
"01001111101010110100111100000011",
"01000111100101000001010001010011",
"00011011110110011000000101001110",
"00101101101001101101101011101100",
"01011100101110110011010101101010",
"01001110000110101100110010000101",
"01011001010101000100001110011101",
"01001100011010010001101111001011",
"01110100101100100001011000011101",
"01011010000101101111101011110101",
"00110100111000000011110100110101",
"00111010001010010110101100011101",
"00001010111011111111010000001010",
"00100101001011110100000100010000",
"01111010110010111110101011010011",
"01011101001000011000111100101110",
"01111001111111000010101100101111",
"01011100101100111010100011011110",
"00101010010100100011011000000001",
"00110100111001111111101001111011",
"01011110111111101001110001010111",
"01001111001101001000011100001000",
"00110010110001001111010110100000",
"00111001000111101100011101110100",
"01001100110110111100010100000000",
"01000110001001111011100010110011",
"00010001010011100101000100101001",
"00101000011001011101000111100000",
"01001000100101011110110111011101",
"01000100000010101000100000000101",
"00000111001010110011110000010100",
"00100011010100010101111011100100",
"01110100110100001011111110011100",
"01011010001000110111011001000000",
"00010011001001110110001000000110",
"00101001010011110000000010100010",
"01000001101110001000101110110001",
"01000000100110011011000110101001",
"00010010110001111001111011000010",
"00101001000111111101100100010101",
"00111010110010010110001110001010",
"00111101001000001000110111111000",
"00010100100110011011101101110010",
"00101010000011000100011011111101",
"00111011101111001100110010000011",
"00111101100110110111010001111010",
"01101101011001010011100010010001",
"01010110011100100011110110011111",
"00000100101100100101111000111001",
"00100010000101110001100110000011",
"01000111101111110110001111001010",
"01000011100111001000010010011101",
"00111111001010110111010010101111",
"00111111010100011000000101111100",
"01101110000110001001001011110100",
"01010110110001011010001000100100",
"01100111100001110100001101000010",
"01010011100000111001010011001101",
"01101110010000101111111001010000",
"01010110110111110110110010001111",
"00111101110000111110000111111000",
"00111110100111100101100000110001",
"00000011011000001100010010010000",
"00100001011011111110000001001010",
"01001010111111100011001110111010",
"01000101001101000110000111101101",
"00010111000110000010010110010101",
"00101011010001010101101101000010",
"01111000000100101101101010101101",
"01011011110000011110010010111001",
"00100010000010000001100110011111",
"00110000101110101010100010111010",
"01110010110111101100010110000001",
"01011001001010001101110011110100",
"01111001110110101001110000011110",
"01011100101001110100011101000100",
"00100001111111010110000000100011",
"00110000101101000001011011001100",
"00011101001100001111101110000010",
"00101110010101001101101100001000",
"01011000110110010011100001110101",
"01001100001001101011111011111001",
"01010100110000100101010111000100",
"01001010000111011011011110111101",
"01101010000011001100000010000010",
"01010100101111011101001010000010",
"01101010001001111000100110011110",
"01010100110011110001100100011011",
"00011101010110000100001110100001",
"00101110011010110100101101110101",
"01110001001101111111110010010110",
"01011000010110010000011011010101",
"01011110111110000100100100111011",
"01001111001100100100010101101100",
"00110000011111111010010110100111",
"00110111111111111101001011001110",
"00110010111100001000100001000111",
"00111001001011110111011100101001",
"01110001101111111110011111111101",
"01011000100111001011101010100001",
"01101011010010010000100100110010",
"01010101011000101101110000000010",
"01000111100010100100001110111010",
"01000011100001010000100010000110",
"00101101011111001011010010000000",
"00110110011111100101100011100010",
"01011000101011100100000111000011",
"01001100000101010101100100100010",
"01001100001111001010000111110011",
"01000101110110111011111111101110",
"01110101001111000001100001001011",
"01011010010110110110111110110001",
"00010111110110011011011001110011",
"00101011101001101110111101001110",
"00111010010101010011010011101000",
"00111100111010011010000000100100",
"01011100110000110101101110001101",
"01001110000111100010000111010011",
"00000110000111001011010011000011",
"00100010110010000100101010101100",
"01111000000110010001011011100000",
"01011011110001011111011110000100",
"01100000001001000010000000011101",
"01001111110011001111101001110010",
"01010001000110101110100001111101",
"01001000010001110010001110101101",
"00001111001100010011110001110101",
"00100111010101010000001000010011",
"01011000001101101111101011001011",
"01001011110110000110111010010100",
"01010000111110010101100101101100",
"01001000001100101010011100001000",
"00110001001110010101011000010100",
"00111000010110011101001000111010",
"01001011000101011100000001001100",
"01000101010000111100101111101011",
"01001010110100111111010110001011",
"01000101001001001011011011010101",
"01010011001101101011011000110111",
"01001001010110000100011000000010",
"01101000010001101011101111001110",
"01010011111000011000111010000001",
"00100011101011010010111000000000",
"00110001100101001110001011000111",
"00100111111110010000101111111011",
"00110011101100101000101101001000",
"01010010010100110111110001010000",
"01001000111010001010111001000010",
"00001101110101001011011110011111",
"00100110101001010000001000101101",
"01000101010100010100111110011101",
"01000010011001110111101100111000",
"01000011100010110111100011100110",
"01000001100001011001110011110000",
"01101100110011010000000011011010",
"01010110001000011111110100101100",
"01110101110100001111010101000100",
"01011010101000111000101101000001",
"01110110011111000000000100101101",
"01011010111111011111111010010011",
"01011110100011001110100011010111",
"01001111000001100100110010111011",
"01100001000110011111111001110110",
"01010000010001101000110100001000",
"00111110000001100100010011100111",
"00111110101110010110011000111000",
"00001100000010011001110101010111",
"00100101101110111011000111011110",
"00111001110010000100000000111010",
"00111100101000000001100110101110",
"00001010010000101110011011011011",
"00100100110111110101111100011110",
"00000001010001011011010110100010",
"00100000011000001111100110000111",
"01010001101000011111011010101101",
"01001000100011111111101111011010",
"01000100100110000001101111000011",
"01000010000010111000100011010101",
"01011110000010010001000100101111",
"01001110101110110101001000110001",
"01010111101111101010101101110000",
"01001011100111000011100100101001",
"00111100101100010011001010100011",
"00111110000101101001101001101001",
"00111110001011010011000101001101",
"00111110110100101001000001110001",
"00101000110110011001001111101101",
"00110100001001101110001000010001",
"01001011111000100110111100011000",
"01000101101010100011111011011011",
"00010110011001000010110000011000",
"00101010111100011010111110011001",
"01111001110100101110110101011001",
"01011100101001000101000000001110",
"01111101000110111100010100101100",
"01011110010001111011000101010011",
"01100001011110011110110001100100",
"01010000011111001111000110000101",
"01000100101001101110001011100100",
"01000010000100100010011111010001",
"01010000010100100111101101100011",
"01000111111010000010000011000001",
"01001001110000001010100000110010",
"01000100100111010000100100001011",
"01101000010101000001000011100101",
"01010011111010001111111111110001",
"01111000010010111000011101011111",
"01011011111001000100001011111001",
"00011100000101000010010010000010",
"00101101110000101011110111111101",
"01110110001010001100100010000100",
"01011010110011111101110111011000",
"00111101100111001101011011111100",
"00111110100011011011000000100000",
"01011111100111111001110101101000",
"01001111100011101110111110011110",
"01100010111101011100100101011110",
"01010001001100010101111100100000",
"00110011011011011100110001000000",
"00111001011101101011101100101010",
"01010110000110111001111010010101",
"01001010110001111001100010010110",
"01000001100000101011001000110101",
"01000000100000010101011101001101",
"00010100100001111100101010110111",
"00101010000000111101011010011111",
"00010100001000011110001101111101",
"00101001110010111001001110100100",
"01001101100011000100111110001100",
"01000110100001100000001110011010",
"01001110010100000000101011110001",
"01000110111001101100011101101011",
"00011110011001001100101001011000",
"00101110111100100000001101011010",
"01001110110100100000010100101111",
"01000111001000111111010110000111",
"00011111111100100000000110011110",
"00101111101100000000000010010110",
"01100010111111001110011000011011",
"01010001001100111110101101101000",
"00101100110110110001011001011110",
"00110110001001110111011000000011",
"01110111101100001010110100001110",
"01011011100101100110000110011010",
"00011111101011100001100010111110",
"00101111100101010100011110001110",
"01101011000010000100011110101011",
"01010101001110101100100001001010",
"00100000100010100100000011111011",
"00110000000001010000011100110100",
"01101011100100001000011111010110",
"01010101100010000000001110101111",
"00000001011011000111001111000011",
"00100000011101100000100000110010",
"00011010010111010010111001010100",
"00101100111011011111010001010111",
"01101000101011000100110100000010",
"01010100000101001000000111110001",
"01100010111001100110000000100111",
"01010001001010111011100010001110",
"01011111000001000001000100111001",
"01001111001101111101111101110010",
"00111000111111101100100001100101",
"00111100001101001001011010100101",
"00101100101001110000100001011001",
"00110110000100100011100000111000",
"01000111010110000010001000011110",
"01000011011010110011100100111001",
"00110001010010100100111111000100",
"00111000011000111001001111111010",
"01001000101110110010110011011011",
"01000100000110101100100011111011",
"00111101100000001110101010100010",
"00111110100000000111010100011011",
"01101110111001110010011011000000",
"01010111001011000000001010000010",
"00101000010110101100101001000011",
"00110011111011001010101000110100",
"00100000011101101011010000000000",
"00101111111110110100111011111111",
"00100010010101001111001100000001",
"00110000111010010111110000000111",
"01111110011101100110100011011001",
"01011110111110110010100010110011",
"01100001111110010110011000110101",
"01010000101100101010101110011101",
"00110110110111001011110110111000",
"00111011001010000001011110000000",
"00010010100110000100110001010110",
"00101001000010111001111100011011",
"00101111100001011011010111000001",
"00110111100000101101001011100111",
"00000101001011001100100010101001",
"00100010010100100101000011001100",
"00110000111111010001011010101110",
"00111000001100111111110010101111",
"01111110010101111011101011110000",
"01011110111010110000000100001101",
"00100101000111101100101001000111",
"00110010010010011001111001111111",
"00010011111110011111110011001001",
"00101001101100101110000110000101",
"00101011001100101101000101001111",
"00110101010101011111010011010000",
"00011100110011110111011101010101",
"00101110001000101111010110000111",
"00110011101010000001010110000111",
"00111001100100101010110111011010",
"00010110001110110001100011111010",
"00101010110110101101101010010000",
"00111101010110011011100001010000",
"00111110011011000001010111011011",
"00011111001110001001110101011101",
"00101111010110010110010110010011",
"00010111101001111000110010111110",
"00101011100100100111001000011111",
"01010111101101101110011010100100",
"01001011100110010000000111110000",
"00000111111001001110101001011111",
"00100011101010110010110100000110",
"01111010100011011110110011100101",
"01011101000001101100100001101111",
"00110110101110101111011111011101",
"00111011000110101011001100010001",
"01000000111000111011001011000100",
"01000000001010101011100001011101",
"00100111001101001111010100111111",
"00110011010101110011101110100101",
"01111110000100110001100111111011",
"01011110110000100000111001111111",
"01110010001011100000001010001001",
"01011000110100110000111101111100",
"01101111111100000010001000011010",
"01010111101011110101000111100001",
"00111011100101000000010010011101",
"00111101100010011010010101000100");

  signal op1,op2,ans1,ans,answ,low,high: std_logic_vector(31 downto 0);
  signal addr: std_logic_vector(19 downto 0) := (others=>'0');
  signal miss: std_logic_vector(31 downto 0) := (others=>'0');
  signal rom_o: std_logic_vector(7 downto 0) := (others=>'1');
  signal uart_go: std_logic;
  signal uart_busy: std_logic := '0';
  signal iter: std_logic_vector(31 downto 0) := (others=>'0');
  signal state: std_logic_vector(4 downto 0) := (others=>'0');
  signal state2: std_logic_vector(4 downto 0) := (others=>'0');

begin

  ib: IBUFG port map (
   i=>MCLK1,
   o=>iclk);
  bg: BUFG port map (
    i=>iclk,
    o=>clk);

  fsqrter:fsqrt port map
    (clk, op1, ans);

  rs232c: u232c generic map (wtime=>x"1ADB")
  port map (
    clk=>clk,
    data=>rom_o,
    go=>uart_go,
    busy=>uart_busy,
    tx=>rs_tx);


 cal: process(clk)
 begin
   if rising_edge(clk) then-- hoge clk後に返答
     if state = "00000" then
       state<=state+1;
       addr<=addr+2;
       op1<=rom(conv_integer(addr));
       ans1<=rom(conv_integer(addr+1));
     elsif state = "00001" then
       state<=state+1;
     elsif state = "00010" then
       state<=state+1;
       answ<=ans;
       state2<="00000";
     elsif state = "00011" and uart_go = '1' then --op1の出力
       state2<=state2+1;
       if op1(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "00100" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "00101" and uart_go = '1' then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "00110" and uart_go = '1' then --op2の出力--nop
       state2<=state2+1;
       if op2(31-conv_integer(state2)) = '1' then
         rom_o<=x"0d";
       else
         rom_o<=x"0d";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "00111" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01000" and uart_go = '1' then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01001" and uart_go = '1' then --outputの出力
       state2<=state2+1;
       if answ(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01010" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01011" and uart_go = '1' then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01100" and uart_go = '1' then --answerの出力
       state2<=state2+1;
       if ans1(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01101" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01110" and uart_go = '1' then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01111" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10000" and uart_go = '1' then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10001" then --low,highとの比較
       state<=state+1;
       low<=ans1 - 3;
     elsif state = "10010" then
       state<=state+1;
       high<=ans1 + 3;
     elsif state = "10011" then
       iter<=iter+1;
       state<=state+1;
       if high < answ or low > answ then
         miss<=miss+1;
       end if;
     elsif state = "10100" and uart_go = '1' then --iterの出力
       state2<=state2+1;
       if iter(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if; 
     elsif state = "10101" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10110" and uart_go = '1' then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10111" and uart_go = '1' then --missの出力
       state2<=state2+1;
       if miss(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "11000" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11001" and uart_go = '1' then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "11010" and uart_go = '1' then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11011" and uart_go = '1' then
       state<="00000";
       rom_o<=x"0a";
     end if;
   end if;
 end process;

    send_msg: process(clk)
  begin
    if rising_edge(clk) then
      if uart_busy='0' and uart_go='0' then
        uart_go<='1';
      else
        uart_go<='0';
      end if;
    end if;
  end process;
  
end VHDL;
