/home/mizuta1018/HW/FPU/VHDL/fsin/fmul_5.vhd