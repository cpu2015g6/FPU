/home/mizuta1018/HW/FPU/VHDL/fsin/revfadd.vhd