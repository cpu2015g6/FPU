/home/mizuta1018/HW/FPU/VHDL/fsin/round1.vhd