library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity invblockram1 is

  generic (
    dwidth : integer := 23;
    awidth : integer := 10);

  port (
    clk  : in  std_logic;
    we   : in  std_logic;
    di   : in  std_logic_vector(dwidth - 1 downto 0);
    do   : out std_logic_vector(dwidth - 1 downto 0);
    addr : in  std_logic_vector(awidth - 1 downto 0));

end invblockram1;

architecture behavioral of invblockram1 is

  type ram_type is
    array(0 to (2 ** awidth) - 1) of std_logic_vector(dwidth - 1 downto 0);

  signal ram : ram_type := ("11111111111111111111110",
"11111111100000000001101",
"11111111000000000111101",
"11111110100000010001101",
"11111110000000011111100",
"11111101100000110001011",
"11111101000001000111001",
"11111100100001100001000",
"11111100000001111110101",
"11111011100010100000001",
"11111011000011000101101",
"11111010100011101111001",
"11111010000100011100010",
"11111001100101001101011",
"11111001000110000010010",
"11111000100110111011001",
"11111000000111110111101",
"11110111101000111000001",
"11110111001001111100100",
"11110110101011000100011",
"11110110001100010000011",
"11110101101101011111111",
"11110101001110110011010",
"11110100110000001010011",
"11110100010001100101010",
"11110011110011000011110",
"11110011010100100110001",
"11110010110110001100001",
"11110010010111110101111",
"11110001111001100011010",
"11110001011011010100011",
"11110000111101001001001",
"11110000011111000001101",
"11110000000000111101101",
"11101111100010111101010",
"11101111000101000000101",
"11101110100111000111100",
"11101110001001010010010",
"11101101101011100000010",
"11101101001101110010000",
"11101100110000000111010",
"11101100010010100000010",
"11101011110100111100110",
"11101011010111011100100",
"11101010111010000000001",
"11101010011100100111001",
"11101001111111010001110",
"11101001100001111111101",
"11101001000100110001010",
"11101000100111100110010",
"11101000001010011110111",
"11100111101101011010111",
"11100111010000011010010",
"11100110110011011101001",
"11100110010110100011100",
"11100101111001101101010",
"11100101011100111010011",
"11100101000000001010111",
"11100100100011011110111",
"11100100000110110110011",
"11100011101010010001001",
"11100011001101101111001",
"11100010110001010000101",
"11100010010100110101100",
"11100001111000011101110",
"11100001011100001001011",
"11100000111111111000000",
"11100000100011101010010",
"11100000000111011111110",
"11011111101011011000101",
"11011111001111010100101",
"11011110110011010011111",
"11011110010111010110100",
"11011101111011011100011",
"11011101011111100101101",
"11011101000011110001111",
"11011100101000000001011",
"11011100001100010100010",
"11011011110000101010011",
"11011011010101000011101",
"11011010111001100000001",
"11011010011101111111101",
"11011010000010100010100",
"11011001100111001000101",
"11011001001011110010000",
"11011000110000011110001",
"11011000010101001101100",
"11010111111010000000010",
"11010111011110110110000",
"11010111000011101110111",
"11010110101000101010111",
"11010110001101101001111",
"11010101110010101100001",
"11010101010111110001011",
"11010100111100111001111",
"11010100100010000101010",
"11010100000111010011101",
"11010011101100100101010",
"11010011010001111010000",
"11010010110111010001101",
"11010010011100101100011",
"11010010000010001001111",
"11010001100111101010101",
"11010001001101001110011",
"11010000110010110101010",
"11010000011000011111000",
"11001111111110001011101",
"11001111100011111011010",
"11001111001001101101111",
"11001110101111100011101",
"11001110010101011100010",
"11001101111011010111110",
"11001101100001010110001",
"11001101000111010111100",
"11001100101101011011111",
"11001100010011100011001",
"11001011111001101101010",
"11001011011111111010011",
"11001011000110001010001",
"11001010101100011101000",
"11001010010010110010110",
"11001001111001001011010",
"11001001011111100110101",
"11001001000110000100110",
"11001000101100100101111",
"11001000010011001010000",
"11000111111001110000110",
"11000111100000011010011",
"11000111000111000110110",
"11000110101101110101111",
"11000110010100101000000",
"11000101111011011100111",
"11000101100010010100100",
"11000101001001001110111",
"11000100110000001100001",
"11000100010111001011111",
"11000011111110001110101",
"11000011100101010100001",
"11000011001100011100011",
"11000010110011100111010",
"11000010011010110101010",
"11000010000010000101010",
"11000001101001011000011",
"11000001010000101110001",
"11000000111000000110101",
"11000000011111100001111",
"11000000000110111111101",
"10111111101110100000010",
"10111111010110000011101",
"10111110111101101001100",
"10111110100101010010001",
"10111110001100111101011",
"10111101110100101011010",
"10111101011100011011101",
"10111101000100001110111",
"10111100101100000100101",
"10111100010011111101001",
"10111011111011111000001",
"10111011100011110110000",
"10111011001011110101111",
"10111010110011111000110",
"10111010011011111110001",
"10111010000100000110001",
"10111001101100010000110",
"10111001010100011101111",
"10111000111100101101100",
"10111000100100111111110",
"10111000001101010100101",
"10110111110101101011111",
"10110111011110000101110",
"10110111000110100010010",
"10110110101111000001000",
"10110110010111100010100",
"10110110000000000110100",
"10110101101000101101000",
"10110101010001010101111",
"10110100111010000001011",
"10110100100010101111010",
"10110100001011011111101",
"10110011110100010010101",
"10110011011101001000000",
"10110011000101111111110",
"10110010101110111010000",
"10110010010111110110110",
"10110010000000110101110",
"10110001101001110111100",
"10110001010010111011100",
"10110000111100000010000",
"10110000100101001010111",
"10110000001110010110001",
"10101111110111100100000",
"10101111100000110011111",
"10101111001010000110011",
"10101110110011011011010",
"10101110011100110010100",
"10101110000110001100001",
"10101101101111101000001",
"10101101011001000110100",
"10101101000010100111010",
"10101100101100001010011",
"10101100010101101111110",
"10101011111111010111100",
"10101011101001000001101",
"10101011010010101110001",
"10101010111100011100111",
"10101010100110001101111",
"10101010010000000001011",
"10101001111001110111000",
"10101001100011101111000",
"10101001001101101001011",
"10101000110111100110000",
"10101000100001100100110",
"10101000001011100110000",
"10100111110101101001011",
"10100111011111101111001",
"10100111001001110111001",
"10100110110100000001011",
"10100110011110001101111",
"10100110001000011100100",
"10100101110010101101100",
"10100101011101000000110",
"10100101000111010110001",
"10100100110001101101110",
"10100100011100000111101",
"10100100000110100011110",
"10100011110001000010001",
"10100011011011100010101",
"10100011000110000101010",
"10100010110000101010010",
"10100010011011010001010",
"10100010000101111010100",
"10100001110000100110001",
"10100001011011010011110",
"10100001000110000011011",
"10100000110000110101011",
"10100000011011101001100",
"10100000000110011111110",
"10011111110001011000001",
"10011111011100010010110",
"10011111000111001111100",
"10011110110010001110010",
"10011110011101001111001",
"10011110001000010010010",
"10011101110011010111100",
"10011101011110011110110",
"10011101001001101000001",
"10011100110100110011110",
"10011100100000000001011",
"10011100001011010001000",
"10011011110110100010110",
"10011011100001110110101",
"10011011001101001100101",
"10011010111000100100101",
"10011010100011111110101",
"10011010001111011010111",
"10011001111010111001011",
"10011001100110011001010",
"10011001010001111011101",
"10011000111101011111111",
"10011000101001000110010",
"10011000010100101110110",
"10011000000000011001001",
"10010111101100000101101",
"10010111010111110100101",
"10010111000011100100101",
"10010110101111010111001",
"10010110011011001011101",
"10010110000111000010010",
"10010101110010111010110",
"10010101011110110101010",
"10010101001010110001111",
"10010100110110110000101",
"10010100100010110000101",
"10010100001110110011001",
"10010011111010110111100",
"10010011100110111101111",
"10010011010011000110001",
"10010010111111010000011",
"10010010101011011100101",
"10010010010111101011001",
"10010010000011111011000",
"10010001110000001101000",
"10010001011100100001000",
"10010001001000110110111",
"10010000110101001110110",
"10010000100001101000100",
"10010000001110000100010",
"10001111111010100001111",
"10001111100111000001001",
"10001111010011100010101",
"10001111000000000101111",
"10001110101100101011001",
"10001110011001010010001",
"10001110000101111011001",
"10001101110010100101111",
"10001101011111010010101",
"10001101001100000001101",
"10001100111000110001101",
"10001100100101100100000",
"10001100010010011000001",
"10001011111111001110001",
"10001011101100000110000",
"10001011011000111111110",
"10001011000101111011011",
"10001010110010111000111",
"10001010011111111000000",
"10001010001100111001000",
"10001001111001111011111",
"10001001100111000000101",
"10001001010100000111001",
"10001001000001001111100",
"10001000101110011001101",
"10001000011011100101101",
"10001000001000110011100",
"10000111110110000010111",
"10000111100011010100010",
"10000111010000100111011",
"10000110111101111100011",
"10000110101011010011000",
"10000110011000101011100",
"10000110000110000101110",
"10000101110011100001111",
"10000101100000111111110",
"10000101001110011111001",
"10000100111100000000011",
"10000100101001100011100",
"10000100010111001000010",
"10000100000100101110111",
"10000011110010010111001",
"10000011100000000001010",
"10000011001101101101000",
"10000010111011011010101",
"10000010101001001001101",
"10000010010110111010101",
"10000010000100101101010",
"10000001110010100001101",
"10000001100000010111110",
"10000001001110001111100",
"10000000111100001001000",
"10000000101010000100011",
"10000000011000000001010",
"10000000000110000000001",
"01111111110100000000000",
"01111111100010000010000",
"01111111010000000101101",
"01111110111110001011000",
"01111110101100010010000",
"01111110011010011010101",
"01111110001000100101000",
"01111101110110110001001",
"01111101100100111110110",
"01111101010011001110000",
"01111101000001011110111",
"01111100101111110001100",
"01111100011110000101110",
"01111100001100011011101",
"01111011111010110011010",
"01111011101001001100011",
"01111011010111100111010",
"01111011000110000011110",
"01111010110100100001111",
"01111010100011000001011",
"01111010010001100010101",
"01111010000000000101100",
"01111001101110101010001",
"01111001011101010000010",
"01111001001011110111111",
"01111000111010100001010",
"01111000101001001100010",
"01111000010111111000110",
"01111000000110100110111",
"01110111110101010110100",
"01110111100100000111110",
"01110111010010111010101",
"01110111000001101111000",
"01110110110000100101000",
"01110110011111011100100",
"01110110001110010101110",
"01110101111101010000011",
"01110101101100001100101",
"01110101011011001010100",
"01110101001010001001110",
"01110100111001001010101",
"01110100101000001101001",
"01110100010111010001001",
"01110100000110010110101",
"01110011110101011101110",
"01110011100100100110010",
"01110011010011110000100",
"01110011000010111100010",
"01110010110010001001011",
"01110010100001011000010",
"01110010010000101000001",
"01110001111111111001111",
"01110001101111001101001",
"01110001011110100001111",
"01110001001101111000001",
"01110000111101001111111",
"01110000101100101001001",
"01110000011100000011110",
"01110000001011100000001",
"01101111111010111101111",
"01101111101010011100111",
"01101111011001111101101",
"01101111001001011111110",
"01101110111001000011011",
"01101110101000101000100",
"01101110011000001111001",
"01101110000111110111001",
"01101101110111100000101",
"01101101100111001011101",
"01101101010110111000000",
"01101101000110100101111",
"01101100110110010101001",
"01101100100110000101111",
"01101100010101111000001",
"01101100000101101011111",
"01101011110101100001000",
"01101011100101010111100",
"01101011010101001111011",
"01101011000101001000111",
"01101010110101000011101",
"01101010100100111111111",
"01101010010100111101100",
"01101010000100111101000",
"01101001110100111101000",
"01101001100100111110111",
"01101001010101000010001",
"01101001000101000111000",
"01101000110101001101001",
"01101000100101010100101",
"01101000010101011101100",
"01101000000101100111111",
"01100111110101110011100",
"01100111100110000000101",
"01100111010110001111001",
"01100111000110011110111",
"01100110110110110000001",
"01100110100111000010110",
"01100110010111010110110",
"01100110000111101100001",
"01100101111000000010111",
"01100101101000011010111",
"01100101011000110100100",
"01100101001001001111011",
"01100100111001101011100",
"01100100101010001001000",
"01100100011010101000001",
"01100100001011001000000",
"01100011111011101001101",
"01100011101100001100100",
"01100011011100110000110",
"01100011001101010110011",
"01100010111101111101010",
"01100010101110100101101",
"01100010011111001111010",
"01100010001111111010001",
"01100010000000100110100",
"01100001110001010100001",
"01100001100010000011001",
"01100001010010110011000",
"01100001000011100100101",
"01100000110100010111011",
"01100000100101001011101",
"01100000010110000001000",
"01100000000110110111110",
"01011111110111101111111",
"01011111101000101001010",
"01011111011001100011111",
"01011111001010011111111",
"01011110111011011101001",
"01011110101100011011101",
"01011110011101011011011",
"01011110001110011100100",
"01011101111111011110111",
"01011101110000100010100",
"01011101100001100111011",
"01011101010010101101101",
"01011101000011110101001",
"01011100110100111101111",
"01011100100110001000000",
"01011100010111010011001",
"01011100001000011111110",
"01011011111001101101100",
"01011011101010111100110",
"01011011011100001100110",
"01011011001101011110010",
"01011010111110110001000",
"01011010110000000101001",
"01011010100001011010011",
"01011010010010110000111",
"01011010000100001000101",
"01011001110101100001101",
"01011001100110111011111",
"01011001011000010111011",
"01011001001001110100000",
"01011000111011010010000",
"01011000101100110001011",
"01011000011110010001010",
"01011000001111110010111",
"01011000000001010101101",
"01010111110010111001101",
"01010111100100011110111",
"01010111010110000101011",
"01010111000111101100111",
"01010110111001010101110",
"01010110101010111111111",
"01010110011100101011000",
"01010110001110010111100",
"01010110000000000101001",
"01010101110001110100000",
"01010101100011100011110",
"01010101010101010101010",
"01010101000111000111110",
"01010100111000111011001",
"01010100101010110000000",
"01010100011100100101110",
"01010100001110011101000",
"01010100000000010101010",
"01010011110010001110101",
"01010011100100001001010",
"01010011010110000101001",
"01010011001000000010000",
"01010010111010000000000",
"01010010101011111111011",
"01010010011101111111110",
"01010010010000000001010",
"01010010000010000100000",
"01010001110100000111111",
"01010001100110001100111",
"01010001011000010011001",
"01010001001010011010100",
"01010000111100100010111",
"01010000101110101100011",
"01010000100000110111010",
"01010000010011000011000",
"01010000000101010000001",
"01001111110111011110001",
"01001111101001101101100",
"01001111011011111101111",
"01001111001110001111011",
"01001111000000100010000",
"01001110110010110101110",
"01001110100101001010101",
"01001110010111100000101",
"01001110001001110111110",
"01001101111100001111111",
"01001101101110101001010",
"01001101100001000011110",
"01001101010011011111010",
"01001101000101111100000",
"01001100111000011001110",
"01001100101010111000100",
"01001100011101011000011",
"01001100001111111001100",
"01001100000010011011101",
"01001011110100111110110",
"01001011100111100011001",
"01001011011010001000100",
"01001011001100101111000",
"01001010111111010110101",
"01001010110001111111010",
"01001010100100101001000",
"01001010010111010011110",
"01001010001001111111101",
"01001001111100101100101",
"01001001101111011010101",
"01001001100010001001110",
"01001001010100111001111",
"01001001000111101011000",
"01001000111010011101011",
"01001000101101010000101",
"01001000100000000101000",
"01001000010010111010100",
"01001000000101110001000",
"01000111111000101000101",
"01000111101011100001010",
"01000111011110011010111",
"01000111010001010101101",
"01000111000100010001011",
"01000110110111001110010",
"01000110101010001100000",
"01000110011101001010111",
"01000110010000001010110",
"01000110000011001011110",
"01000101110110001101110",
"01000101101001010000101",
"01000101011100010100110",
"01000101001111011001110",
"01000101000010011111111",
"01000100110101100111000",
"01000100101000101111010",
"01000100011011111000011",
"01000100001111000010100",
"01000100000010001101110",
"01000011110101011010000",
"01000011101000100111010",
"01000011011011110101011",
"01000011001111000100101",
"01000011000010010100111",
"01000010110101100110001",
"01000010101000111000010",
"01000010011100001011100",
"01000010001111011111111",
"01000010000010110101001",
"01000001110110001011011",
"01000001101001100010101",
"01000001011100111010110",
"01000001010000010100000",
"01000001000011101110010",
"01000000110111001001100",
"01000000101010100101101",
"01000000011110000010110",
"01000000010001100000111",
"01000000000101000000001",
"00111111111000100000000",
"00111111101100000001001",
"00111111011111100011001",
"00111111010011000110001",
"00111111000110101010010",
"00111110111010001111001",
"00111110101101110101001",
"00111110100001011100000",
"00111110010101000011111",
"00111110001000101100101",
"00111101111100010110100",
"00111101110000000001010",
"00111101100011101100111",
"00111101010111011001101",
"00111101001011000111001",
"00111100111110110101101",
"00111100110010100101010",
"00111100100110010101100",
"00111100011010000110111",
"00111100001101111001010",
"00111100000001101100100",
"00111011110101100000110",
"00111011101001010101111",
"00111011011101001100000",
"00111011010001000011001",
"00111011000100111011000",
"00111010111000110011111",
"00111010101100101101110",
"00111010100000101000100",
"00111010010100100100001",
"00111010001000100000110",
"00111001111100011110011",
"00111001110000011100110",
"00111001100100011100010",
"00111001011000011100011",
"00111001001100011101100",
"00111001000000011111101",
"00111000110100100010110",
"00111000101000100110101",
"00111000011100101011100",
"00111000010000110001011",
"00111000000100110111111",
"00110111111000111111101",
"00110111101101001000001",
"00110111100001010001100",
"00110111010101011011110",
"00110111001001100110111",
"00110110111101110011000",
"00110110110010000000000",
"00110110100110001101111",
"00110110011010011100101",
"00110110001110101100001",
"00110110000010111100111",
"00110101110111001110010",
"00110101101011100000100",
"00110101011111110011110",
"00110101010100000111111",
"00110101001000011100111",
"00110100111100110010110",
"00110100110001001001100",
"00110100100101100001001",
"00110100011001111001101",
"00110100001110010011000",
"00110100000010101101010",
"00110011110111001000010",
"00110011101011100100010",
"00110011100000000001001",
"00110011010100011110110",
"00110011001000111101011",
"00110010111101011101000",
"00110010110001111101001",
"00110010100110011110010",
"00110010011011000000010",
"00110010001111100011001",
"00110010000100000110111",
"00110001111000101011100",
"00110001101101010001000",
"00110001100001110111010",
"00110001010110011110011",
"00110001001011000110011",
"00110000111111101111010",
"00110000110100011001000",
"00110000101001000011100",
"00110000011101101110110",
"00110000010010011011000",
"00110000000111001000001",
"00101111111011110110000",
"00101111110000100100101",
"00101111100101010100011",
"00101111011010000100100",
"00101111001110110101110",
"00101111000011100111111",
"00101110111000011010110",
"00101110101101001110100",
"00101110100010000011000",
"00101110010110111000011",
"00101110001011101110101",
"00101110000000100101101",
"00101101110101011101100",
"00101101101010010110010",
"00101101011111001111100",
"00101101010100001010000",
"00101101001001000101000",
"00101100111110000001000",
"00101100110010111101101",
"00101100100111111011010",
"00101100011100111001100",
"00101100010001111000110",
"00101100000110111000101",
"00101011111011111001011",
"00101011110000111011000",
"00101011100101111101011",
"00101011011011000000100",
"00101011010000000100100",
"00101011000101001001011",
"00101010111010001110111",
"00101010101111010101010",
"00101010100100011100011",
"00101010011001100100100",
"00101010001110101101001",
"00101010000011110110110",
"00101001111001000001001",
"00101001101110001100001",
"00101001100011011000001",
"00101001011000100100110",
"00101001001101110010011",
"00101001000011000000100",
"00101000111000001111100",
"00101000101101011111011",
"00101000100010110000000",
"00101000011000000001010",
"00101000001101010011100",
"00101000000010100110011",
"00100111110111111010001",
"00100111101101001110101",
"00100111100010100011110",
"00100111010111111001110",
"00100111001101010000100",
"00100111000010101000010",
"00100110111000000000100",
"00100110101101011001100",
"00100110100010110011011",
"00100110011000001110000",
"00100110001101101001011",
"00100110000011000101100",
"00100101111000100010010",
"00100101101110000000000",
"00100101100011011110011",
"00100101011000111101100",
"00100101001110011101010",
"00100101000011111110000",
"00100100111001011111011",
"00100100101111000001100",
"00100100100100100100011",
"00100100011010001000001",
"00100100001111101100011",
"00100100000101010001101",
"00100011111010110111100",
"00100011110000011110001",
"00100011100110000101011",
"00100011011011101101101",
"00100011010001010110011",
"00100011000110111111111",
"00100010111100101010010",
"00100010110010010101010",
"00100010101000000001000",
"00100010011101101101101",
"00100010010011011010110",
"00100010001001001000110",
"00100001111110110111011",
"00100001110100100110111",
"00100001101010010110111",
"00100001100000000111110",
"00100001010101111001011",
"00100001001011101011101",
"00100001000001011110101",
"00100000110111010010100",
"00100000101101000110111",
"00100000100010111100001",
"00100000011000110010000",
"00100000001110101000101",
"00100000000100011111111",
"00011111111010011000000",
"00011111110000010000110",
"00011111100110001010010",
"00011111011100000100011",
"00011111010001111111010",
"00011111000111111010111",
"00011110111101110111001",
"00011110110011110100001",
"00011110101001110001111",
"00011110011111110000010",
"00011110010101101111010",
"00011110001011101111000",
"00011110000001101111100",
"00011101110111110000110",
"00011101101101110010101",
"00011101100011110101010",
"00011101011001111000100",
"00011101001111111100100",
"00011101000110000001001",
"00011100111100000110100",
"00011100110010001100100",
"00011100101000010011010",
"00011100011110011010110",
"00011100010100100010111",
"00011100001010101011101",
"00011100000000110101001",
"00011011110110111111010",
"00011011101101001010001",
"00011011100011010101101",
"00011011011001100001111",
"00011011001111101110110",
"00011011000101111100010",
"00011010111100001010100",
"00011010110010011001100",
"00011010101000101001001",
"00011010011110111001001",
"00011010010101001010001",
"00011010001011011011110",
"00011010000001101110000",
"00011001111000000000111",
"00011001101110010100101",
"00011001100100101000111",
"00011001011010111101110",
"00011001010001010011011",
"00011001000111101001101",
"00011000111110000000100",
"00011000110100011000001",
"00011000101010110000011",
"00011000100001001001010",
"00011000010111100010110",
"00011000001101111101001",
"00011000000100010111111",
"00010111111010110011100",
"00010111110001001111101",
"00010111100111101100100",
"00010111011110001010000",
"00010111010100101000001",
"00010111001011000110111",
"00010111000001100110011",
"00010110111000000110011",
"00010110101110100111000",
"00010110100101001000100",
"00010110011011101010100",
"00010110010010001101001",
"00010110001000110000100",
"00010101111111010100011",
"00010101110101111000111",
"00010101101100011110001",
"00010101100011000100000",
"00010101011001101010100",
"00010101010000010001101",
"00010101000110111001100",
"00010100111101100001111",
"00010100110100001011000",
"00010100101010110100101",
"00010100100001011111000",
"00010100011000001001111",
"00010100001110110101011",
"00010100000101100001101",
"00010011111100001110011",
"00010011110010111011111",
"00010011101001101001111",
"00010011100000011000101",
"00010011010111001000000",
"00010011001101110111110",
"00010011000100101000011",
"00010010111011011001101",
"00010010110010001011011",
"00010010101000111101110",
"00010010011111110000111",
"00010010010110100100100",
"00010010001101011000110",
"00010010000100001101101",
"00010001111011000011001",
"00010001110001111001001",
"00010001101000101111111",
"00010001011111100111010",
"00010001010110011111010",
"00010001001101010111110",
"00010001000100010000111",
"00010000111011001010101",
"00010000110010000101000",
"00010000101001000000000",
"00010000011111111011101",
"00010000010110110111110",
"00010000001101110100100",
"00010000000100110010000",
"00001111111011110000000",
"00001111110010101110100",
"00001111101001101101101",
"00001111100000101101011",
"00001111010111101101110",
"00001111001110101110110",
"00001111000101110000011",
"00001110111100110010100",
"00001110110011110101010",
"00001110101010111000100",
"00001110100001111100100",
"00001110011001000001000",
"00001110010000000110001",
"00001110000111001011111",
"00001101111110010010001",
"00001101110101011001000",
"00001101101100100000100",
"00001101100011101000101",
"00001101011010110001001",
"00001101010001111010011",
"00001101001001000100001",
"00001101000000001110100",
"00001100110111011001100",
"00001100101110100101000",
"00001100100101110001001",
"00001100011100111101111",
"00001100010100001011001",
"00001100001011011001000",
"00001100000010100111011",
"00001011111001110110011",
"00001011110001000110001",
"00001011101000010110000",
"00001011011111100110110",
"00001011010110111000000",
"00001011001110001001110",
"00001011000101011100010",
"00001010111100101111010",
"00001010110100000010110",
"00001010101011010110111",
"00001010100010101011101",
"00001010011010000000110",
"00001010010001010110101",
"00001010001000101101000",
"00001010000000000100000",
"00001001110111011011100",
"00001001101110110011100",
"00001001100110001100001",
"00001001011101100101011",
"00001001010100111111000",
"00001001001100011001011",
"00001001000011110100010",
"00001000111011001111101",
"00001000110010101011100",
"00001000101010001000000",
"00001000100001100101001",
"00001000011001000010110",
"00001000010000100000111",
"00001000000111111111101",
"00000111111111011110111",
"00000111110110111110100",
"00000111101110011110111",
"00000111100101111111111",
"00000111011101100001011",
"00000111010101000011010",
"00000111001100100101111",
"00000111000100001000111",
"00000110111011101100100",
"00000110110011010000101",
"00000110101010110101011",
"00000110100010011010101",
"00000110011010000000011",
"00000110010001100110110",
"00000110001001001101101",
"00000110000000110101000",
"00000101111000011101000",
"00000101110000000101100",
"00000101100111101110011",
"00000101011111011000000",
"00000101010111000010000",
"00000101001110101100101",
"00000101000110010111110",
"00000100111110000011100",
"00000100110101101111101",
"00000100101101011100011",
"00000100100101001001101",
"00000100011100110111011",
"00000100010100100101110",
"00000100001100010100101",
"00000100000100000100000",
"00000011111011110011110",
"00000011110011100100001",
"00000011101011010101001",
"00000011100011000110100",
"00000011011010111000100",
"00000011010010101011000",
"00000011001010011101111",
"00000011000010010001100",
"00000010111010000101100",
"00000010110001111010001",
"00000010101001101111001",
"00000010100001100100110",
"00000010011001011010111",
"00000010010001010001100",
"00000010001001001000101",
"00000010000001000000011",
"00000001111000111000100",
"00000001110000110001001",
"00000001101000101010011",
"00000001100000100100001",
"00000001011000011110010",
"00000001010000011001000",
"00000001001000010100010",
"00000001000000010000000",
"00000000111000001100001",
"00000000110000001000111",
"00000000101000000110001",
"00000000100000000100000",
"00000000011000000010001",
"00000000010000000000111",
"00000000001000000000001");

  signal reg_addr : std_logic_vector(awidth - 1 downto 0);

begin

  process(clk)
  begin
    if rising_edge(clk) then
      if we = '1' then
        ram(conv_integer(addr)) <= di;
      end if;
      reg_addr <= addr;
    end if;
  end process;

  do <= ram(conv_integer(reg_addr));

end behavioral;
