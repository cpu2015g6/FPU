/home/mizuta1018/HW/FPU/VHDL/finv/fmul_inv.vhd