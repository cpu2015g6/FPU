/home/mizuta1018/HW/FPU/VHDL/finv/quamul.vhd