/home/mizuta1018/HW/FPU/VHDL/fsin/kernel_cos.vhd