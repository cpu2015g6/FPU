/home/mizuta1018/HW/FPU/VHDL/fsin/round2.vhd