/home/mizuta1018/HW/FPU/VHDL/fcos/fadd.vhd