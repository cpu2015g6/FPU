library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

entity sqrtromfetch is
  port(addr: in std_logic_vector(10 downto 0);
       data,data2:  out std_logic_vector(22 downto 0) -- 23bit
       );
  end sqrtromfetch;

architecture VHDL of sqrtromfetch is

  type rom_t is array(0 to 2047) of std_logic_vector(22 downto 0);
  constant rom1 : rom_t :=("00000000000000000000000",
"00000000000111111111111",
"00000000001111111111100",
"00000000010111111110111",
"00000000011111111110000",
"00000000100111111100111",
"00000000101111111011100",
"00000000110111111001111",
"00000000111111111000000",
"00000001000111110101111",
"00000001001111110011100",
"00000001010111110000111",
"00000001011111101110001",
"00000001100111101011000",
"00000001101111100111101",
"00000001110111100100000",
"00000001111111100000010",
"00000010000111011100001",
"00000010001111010111111",
"00000010010111010011010",
"00000010011111001110100",
"00000010100111001001011",
"00000010101111000100001",
"00000010110110111110101",
"00000010111110111000110",
"00000011000110110010110",
"00000011001110101100100",
"00000011010110100110000",
"00000011011110011111010",
"00000011100110011000010",
"00000011101110010001001",
"00000011110110001001101",
"00000011111110000001111",
"00000100000101111010000",
"00000100001101110001111",
"00000100010101101001011",
"00000100011101100000110",
"00000100100101010111111",
"00000100101101001110110",
"00000100110101000101011",
"00000100111100111011110",
"00000101000100110010000",
"00000101001100100111111",
"00000101010100011101101",
"00000101011100010011000",
"00000101100100001000010",
"00000101101011111101010",
"00000101110011110010000",
"00000101111011100110100",
"00000110000011011010111",
"00000110001011001110111",
"00000110010011000010110",
"00000110011010110110010",
"00000110100010101001101",
"00000110101010011100110",
"00000110110010001111101",
"00000110111010000010011",
"00000111000001110100110",
"00000111001001100111000",
"00000111010001011001000",
"00000111011001001010110",
"00000111100000111100010",
"00000111101000101101100",
"00000111110000011110100",
"00000111111000001111011",
"00001000000000000000000",
"00001000000111110000011",
"00001000001111100000100",
"00001000010111010000011",
"00001000011111000000001",
"00001000100110101111100",
"00001000101110011110110",
"00001000110110001101110",
"00001000111101111100101",
"00001001000101101011001",
"00001001001101011001100",
"00001001010101000111101",
"00001001011100110101100",
"00001001100100100011001",
"00001001101100010000100",
"00001001110011111101110",
"00001001111011101010110",
"00001010000011010111100",
"00001010001011000100001",
"00001010010010110000011",
"00001010011010011100100",
"00001010100010001000011",
"00001010101001110100000",
"00001010110001011111100",
"00001010111001001010101",
"00001011000000110101101",
"00001011001000100000011",
"00001011010000001011000",
"00001011010111110101011",
"00001011011111011111011",
"00001011100111001001011",
"00001011101110110011000",
"00001011110110011100100",
"00001011111110000101110",
"00001100000101101110110",
"00001100001101010111100",
"00001100010101000000001",
"00001100011100101000100",
"00001100100100010000101",
"00001100101011111000100",
"00001100110011100000010",
"00001100111011000111110",
"00001101000010101111000",
"00001101001010010110001",
"00001101010001111101000",
"00001101011001100011101",
"00001101100001001010000",
"00001101101000110000010",
"00001101110000010110010",
"00001101110111111100000",
"00001101111111100001101",
"00001110000111000111000",
"00001110001110101100001",
"00001110010110010001001",
"00001110011101110101110",
"00001110100101011010010",
"00001110101100111110101",
"00001110110100100010101",
"00001110111100000110100",
"00001111000011101010010",
"00001111001011001101101",
"00001111010010110000111",
"00001111011010010100000",
"00001111100001110110110",
"00001111101001011001011",
"00001111110000111011110",
"00001111111000011110000",
"00010000000000000000000",
"00010000000111100001110",
"00010000001111000011011",
"00010000010110100100101",
"00010000011110000101111",
"00010000100101100110110",
"00010000101101000111100",
"00010000110100101000000",
"00010000111100001000011",
"00010001000011101000100",
"00010001001011001000011",
"00010001010010101000001",
"00010001011010000111101",
"00010001100001100110111",
"00010001101001000110000",
"00010001110000100100111",
"00010001111000000011101",
"00010001111111100010001",
"00010010000111000000011",
"00010010001110011110011",
"00010010010101111100010",
"00010010011101011010000",
"00010010100100110111011",
"00010010101100010100101",
"00010010110011110001110",
"00010010111011001110101",
"00010011000010101011010",
"00010011001010000111110",
"00010011010001100100000",
"00010011011001000000000",
"00010011100000011011111",
"00010011100111110111100",
"00010011101111010011000",
"00010011110110101110001",
"00010011111110001001010",
"00010100000101100100001",
"00010100001100111110110",
"00010100010100011001001",
"00010100011011110011011",
"00010100100011001101100",
"00010100101010100111011",
"00010100110010000001000",
"00010100111001011010100",
"00010101000000110011110",
"00010101001000001100110",
"00010101001111100101101",
"00010101010110111110011",
"00010101011110010110110",
"00010101100101101111001",
"00010101101101000111001",
"00010101110100011111000",
"00010101111011110110110",
"00010110000011001110010",
"00010110001010100101100",
"00010110010001111100101",
"00010110011001010011100",
"00010110100000101010010",
"00010110101000000000110",
"00010110101111010111001",
"00010110110110101101010",
"00010110111110000011001",
"00010111000101011000111",
"00010111001100101110100",
"00010111010100000011111",
"00010111011011011001000",
"00010111100010101110000",
"00010111101010000010110",
"00010111110001010111011",
"00010111111000101011110",
"00011000000000000000000",
"00011000000111010100000",
"00011000001110100111111",
"00011000010101111011100",
"00011000011101001110111",
"00011000100100100010001",
"00011000101011110101010",
"00011000110011001000001",
"00011000111010011010110",
"00011001000001101101010",
"00011001001000111111101",
"00011001010000010001110",
"00011001010111100011101",
"00011001011110110101011",
"00011001100110000111000",
"00011001101101011000011",
"00011001110100101001100",
"00011001111011111010100",
"00011010000011001011010",
"00011010001010011011111",
"00011010010001101100011",
"00011010011000111100101",
"00011010100000001100101",
"00011010100111011100100",
"00011010101110101100010",
"00011010110101111011110",
"00011010111101001011000",
"00011011000100011010001",
"00011011001011101001001",
"00011011010010110111111",
"00011011011010000110100",
"00011011100001010100111",
"00011011101000100011000",
"00011011101111110001001",
"00011011110110111110111",
"00011011111110001100101",
"00011100000101011010000",
"00011100001100100111011",
"00011100010011110100100",
"00011100011011000001011",
"00011100100010001110001",
"00011100101001011010110",
"00011100110000100111001",
"00011100110111110011010",
"00011100111110111111010",
"00011101000110001011001",
"00011101001101010110110",
"00011101010100100010010",
"00011101011011101101100",
"00011101100010111000101",
"00011101101010000011101",
"00011101110001001110011",
"00011101111000011000111",
"00011101111111100011011",
"00011110000110101101100",
"00011110001101110111101",
"00011110010101000001011",
"00011110011100001011001",
"00011110100011010100101",
"00011110101010011101111",
"00011110110001100111001",
"00011110111000110000000",
"00011110111111111000111",
"00011111000111000001100",
"00011111001110001001111",
"00011111010101010010001",
"00011111011100011010010",
"00011111100011100010001",
"00011111101010101001111",
"00011111110001110001011",
"00011111111000111000110",
"00100000000000000000000",
"00100000000111000111000",
"00100000001110001101111",
"00100000010101010100100",
"00100000011100011011000",
"00100000100011100001011",
"00100000101010100111100",
"00100000110001101101100",
"00100000111000110011010",
"00100000111111111000111",
"00100001000110111110011",
"00100001001110000011101",
"00100001010101001000110",
"00100001011100001101101",
"00100001100011010010011",
"00100001101010010111000",
"00100001110001011011011",
"00100001111000011111101",
"00100001111111100011110",
"00100010000110100111101",
"00100010001101101011011",
"00100010010100101110111",
"00100010011011110010010",
"00100010100010110101100",
"00100010101001111000100",
"00100010110000111011011",
"00100010110111111110001",
"00100010111111000000101",
"00100011000110000011000",
"00100011001101000101001",
"00100011010100000111001",
"00100011011011001001000",
"00100011100010001010110",
"00100011101001001100010",
"00100011110000001101101",
"00100011110111001110110",
"00100011111110001111110",
"00100100000101010000101",
"00100100001100010001010",
"00100100010011010001110",
"00100100011010010010001",
"00100100100001010010010",
"00100100101000010010010",
"00100100101111010010000",
"00100100110110010001110",
"00100100111101010001010",
"00100101000100010000100",
"00100101001011001111110",
"00100101010010001110110",
"00100101011001001101100",
"00100101100000001100001",
"00100101100111001010101",
"00100101101110001001000",
"00100101110101000111001",
"00100101111100000101001",
"00100110000011000011000",
"00100110001010000000101",
"00100110010000111110001",
"00100110010111111011100",
"00100110011110111000101",
"00100110100101110101110",
"00100110101100110010100",
"00100110110011101111010",
"00100110111010101011110",
"00100111000001101000001",
"00100111001000100100010",
"00100111001111100000011",
"00100111010110011100001",
"00100111011101010111111",
"00100111100100010011011",
"00100111101011001110110",
"00100111110010001010000",
"00100111111001000101001",
"00101000000000000000000",
"00101000000110111010110",
"00101000001101110101010",
"00101000010100101111101",
"00101000011011101001111",
"00101000100010100100000",
"00101000101001011101111",
"00101000110000010111110",
"00101000110111010001010",
"00101000111110001010110",
"00101001000101000100000",
"00101001001011111101001",
"00101001010010110110001",
"00101001011001101110111",
"00101001100000100111100",
"00101001100111100000000",
"00101001101110011000011",
"00101001110101010000100",
"00101001111100001000100",
"00101010000011000000011",
"00101010001001111000001",
"00101010010000101111101",
"00101010010111100111000",
"00101010011110011110010",
"00101010100101010101010",
"00101010101100001100001",
"00101010110011000010111",
"00101010111001111001100",
"00101011000000101111111",
"00101011000111100110001",
"00101011001110011100010",
"00101011010101010010010",
"00101011011100001000000",
"00101011100010111101110",
"00101011101001110011010",
"00101011110000101000100",
"00101011110111011101110",
"00101011111110010010110",
"00101100000101000111101",
"00101100001011111100011",
"00101100010010110000111",
"00101100011001100101010",
"00101100100000011001100",
"00101100100111001101101",
"00101100101110000001100",
"00101100110100110101011",
"00101100111011101001000",
"00101101000010011100100",
"00101101001001001111110",
"00101101010000000011000",
"00101101010110110110000",
"00101101011101101000111",
"00101101100100011011100",
"00101101101011001110001",
"00101101110010000000100",
"00101101111000110010110",
"00101101111111100100111",
"00101110000110010110110",
"00101110001101001000101",
"00101110010011111010010",
"00101110011010101011110",
"00101110100001011101000",
"00101110101000001110010",
"00101110101110111111010",
"00101110110101110000001",
"00101110111100100000111",
"00101111000011010001100",
"00101111001010000001111",
"00101111010000110010010",
"00101111010111100010011",
"00101111011110010010010",
"00101111100101000010001",
"00101111101011110001111",
"00101111110010100001011",
"00101111111001010000110",
"00110000000000000000000",
"00110000000110101111000",
"00110000001101011110000",
"00110000010100001100110",
"00110000011010111011011",
"00110000100001101001111",
"00110000101000011000010",
"00110000101111000110011",
"00110000110101110100100",
"00110000111100100010011",
"00110001000011010000001",
"00110001001001111101110",
"00110001010000101011001",
"00110001010111011000100",
"00110001011110000101101",
"00110001100100110010101",
"00110001101011011111100",
"00110001110010001100010",
"00110001111000111000110",
"00110001111111100101010",
"00110010000110010001100",
"00110010001100111101101",
"00110010010011101001101",
"00110010011010010101011",
"00110010100001000001001",
"00110010100111101100101",
"00110010101110011000000",
"00110010110101000011010",
"00110010111011101110011",
"00110011000010011001011",
"00110011001001000100010",
"00110011001111101110111",
"00110011010110011001011",
"00110011011101000011110",
"00110011100011101110000",
"00110011101010011000001",
"00110011110001000010001",
"00110011110111101011111",
"00110011111110010101101",
"00110100000100111111001",
"00110100001011101000100",
"00110100010010010001110",
"00110100011000111010110",
"00110100011111100011110",
"00110100100110001100100",
"00110100101100110101010",
"00110100110011011101110",
"00110100111010000110001",
"00110101000000101110011",
"00110101000111010110100",
"00110101001101111110011",
"00110101010100100110010",
"00110101011011001101111",
"00110101100001110101011",
"00110101101000011100110",
"00110101101111000100000",
"00110101110101101011001",
"00110101111100010010001",
"00110110000010111000111",
"00110110001001011111101",
"00110110010000000110001",
"00110110010110101100100",
"00110110011101010010110",
"00110110100011111000111",
"00110110101010011110111",
"00110110110001000100110",
"00110110110111101010100",
"00110110111110010000000",
"00110111000100110101011",
"00110111001011011010110",
"00110111010001111111111",
"00110111011000100100111",
"00110111011111001001110",
"00110111100101101110100",
"00110111101100010011000",
"00110111110010110111100",
"00110111111001011011110",
"00111000000000000000000",
"00111000000110100100000",
"00111000001101000111111",
"00111000010011101011101",
"00111000011010001111010",
"00111000100000110010110",
"00111000100111010110001",
"00111000101101111001010",
"00111000110100011100011",
"00111000111010111111010",
"00111001000001100010001",
"00111001001000000100110",
"00111001001110100111010",
"00111001010101001001101",
"00111001011011101011111",
"00111001100010001110000",
"00111001101000110000000",
"00111001101111010001111",
"00111001110101110011101",
"00111001111100010101001",
"00111010000010110110101",
"00111010001001010111111",
"00111010001111111001000",
"00111010010110011010001",
"00111010011100111011000",
"00111010100011011011110",
"00111010101001111100011",
"00111010110000011100111",
"00111010110110111101010",
"00111010111101011101011",
"00111011000011111101100",
"00111011001010011101100",
"00111011010000111101010",
"00111011010111011101000",
"00111011011101111100100",
"00111011100100011011111",
"00111011101010111011010",
"00111011110001011010011",
"00111011110111111001011",
"00111011111110011000010",
"00111100000100110111000",
"00111100001011010101101",
"00111100010001110100001",
"00111100011000010010100",
"00111100011110110000110",
"00111100100101001110110",
"00111100101011101100110",
"00111100110010001010101",
"00111100111000101000010",
"00111100111111000101111",
"00111101000101100011010",
"00111101001100000000100",
"00111101010010011101110",
"00111101011000111010110",
"00111101011111010111101",
"00111101100101110100011",
"00111101101100010001000",
"00111101110010101101101",
"00111101111001001010000",
"00111101111111100110010",
"00111110000110000010011",
"00111110001100011110010",
"00111110010010111010001",
"00111110011001010101111",
"00111110011111110001100",
"00111110100110001101000",
"00111110101100101000010",
"00111110110011000011100",
"00111110111001011110101",
"00111110111111111001100",
"00111111000110010100011",
"00111111001100101111000",
"00111111010011001001101",
"00111111011001100100000",
"00111111011111111110011",
"00111111100110011000100",
"00111111101100110010101",
"00111111110011001100100",
"00111111111001100110010",
"01000000000000000000000",
"01000000000110011001100",
"01000000001100110010111",
"01000000010011001100001",
"01000000011001100101011",
"01000000011111111110011",
"01000000100110010111010",
"01000000101100110000000",
"01000000110011001000101",
"01000000111001100001010",
"01000000111111111001101",
"01000001000110010001111",
"01000001001100101010000",
"01000001010011000010000",
"01000001011001011001111",
"01000001011111110001101",
"01000001100110001001010",
"01000001101100100000110",
"01000001110010111000001",
"01000001111001001111011",
"01000001111111100110100",
"01000010000101111101100",
"01000010001100010100011",
"01000010010010101011001",
"01000010011001000001110",
"01000010011111011000010",
"01000010100101101110101",
"01000010101100000100111",
"01000010110010011011000",
"01000010111000110001000",
"01000010111111000110111",
"01000011000101011100101",
"01000011001011110010010",
"01000011010010000111110",
"01000011011000011101001",
"01000011011110110010011",
"01000011100101000111100",
"01000011101011011100100",
"01000011110001110001011",
"01000011111000000110001",
"01000011111110011010111",
"01000100000100101111011",
"01000100001011000011110",
"01000100010001011000000",
"01000100010111101100001",
"01000100011110000000001",
"01000100100100010100000",
"01000100101010100111111",
"01000100110000111011100",
"01000100110111001111000",
"01000100111101100010011",
"01000101000011110101110",
"01000101001010001000111",
"01000101010000011011111",
"01000101010110101110111",
"01000101011101000001101",
"01000101100011010100010",
"01000101101001100110111",
"01000101101111111001010",
"01000101110110001011101",
"01000101111100011101110",
"01000110000010101111111",
"01000110001001000001110",
"01000110001111010011101",
"01000110010101100101011",
"01000110011011110110111",
"01000110100010001000011",
"01000110101000011001110",
"01000110101110101011000",
"01000110110100111100000",
"01000110111011001101000",
"01000111000001011101111",
"01000111000111101110101",
"01000111001101111111010",
"01000111010100001111110",
"01000111011010100000001",
"01000111100000110000011",
"01000111100111000000101",
"01000111101101010000101",
"01000111110011100000100",
"01000111111001110000010",
"01001000000000000000000",
"01001000000110001111100",
"01001000001100011111000",
"01001000010010101110010",
"01001000011000111101100",
"01001000011111001100100",
"01001000100101011011100",
"01001000101011101010011",
"01001000110001111001000",
"01001000111000000111101",
"01001000111110010110001",
"01001001000100100100100",
"01001001001010110010110",
"01001001010001000000111",
"01001001010111001110111",
"01001001011101011100110",
"01001001100011101010101",
"01001001101001111000010",
"01001001110000000101110",
"01001001110110010011010",
"01001001111100100000100",
"01001010000010101101110",
"01001010001000111010110",
"01001010001111000111110",
"01001010010101010100101",
"01001010011011100001011",
"01001010100001101110000",
"01001010100111111010100",
"01001010101110000110111",
"01001010110100010011001",
"01001010111010011111010",
"01001011000000101011010",
"01001011000110110111010",
"01001011001101000011000",
"01001011010011001110101",
"01001011011001011010010",
"01001011011111100101110",
"01001011100101110001000",
"01001011101011111100010",
"01001011110010000111011",
"01001011111000010010011",
"01001011111110011101010",
"01001100000100101000000",
"01001100001010110010101",
"01001100010000111101010",
"01001100010111000111101",
"01001100011101010010000",
"01001100100011011100001",
"01001100101001100110010",
"01001100101111110000010",
"01001100110101111010000",
"01001100111100000011110",
"01001101000010001101011",
"01001101001000010110111",
"01001101001110100000011",
"01001101010100101001101",
"01001101011010110010110",
"01001101100000111011111",
"01001101100111000100110",
"01001101101101001101101",
"01001101110011010110011",
"01001101111001011111000",
"01001101111111100111011",
"01001110000101101111111",
"01001110001011111000001",
"01001110010010000000010",
"01001110011000001000010",
"01001110011110010000010",
"01001110100100011000000",
"01001110101010011111110",
"01001110110000100111011",
"01001110110110101110111",
"01001110111100110110010",
"01001111000010111101100",
"01001111001001000100101",
"01001111001111001011101",
"01001111010101010010101",
"01001111011011011001011",
"01001111100001100000001",
"01001111100111100110110",
"01001111101101101101001",
"01001111110011110011100",
"01001111111001111001110",
"01010000000000000000000",
"01010000000110000110000",
"01010000001100001011111",
"01010000010010010001110",
"01010000011000010111100",
"01010000011110011101000",
"01010000100100100010100",
"01010000101010100111111",
"01010000110000101101010",
"01010000110110110010011",
"01010000111100110111011",
"01010001000010111100011",
"01010001001001000001001",
"01010001001111000101111",
"01010001010101001010100",
"01010001011011001111000",
"01010001100001010011011",
"01010001100111010111101",
"01010001101101011011111",
"01010001110011011111111",
"01010001111001100011111",
"01010001111111100111110",
"01010010000101101011100",
"01010010001011101111001",
"01010010010001110010101",
"01010010010111110110000",
"01010010011101111001011",
"01010010100011111100100",
"01010010101001111111101",
"01010010110000000010101",
"01010010110110000101100",
"01010010111100001000010",
"01010011000010001010111",
"01010011001000001101100",
"01010011001110001111111",
"01010011010100010010010",
"01010011011010010100100",
"01010011100000010110101",
"01010011100110011000101",
"01010011101100011010100",
"01010011110010011100010",
"01010011111000011110000",
"01010011111110011111101",
"01010100000100100001000",
"01010100001010100010011",
"01010100010000100011110",
"01010100010110100100111",
"01010100011100100101111",
"01010100100010100110111",
"01010100101000100111110",
"01010100101110101000011",
"01010100110100101001000",
"01010100111010101001101",
"01010101000000101010000",
"01010101000110101010010",
"01010101001100101010100",
"01010101010010101010101",
"01010101011000101010101",
"01010101011110101010100",
"01010101100100101010010",
"01010101101010101010000",
"01010101110000101001100",
"01010101110110101001000",
"01010101111100101000011",
"01010110000010100111101",
"01010110001000100110110",
"01010110001110100101111",
"01010110010100100100110",
"01010110011010100011101",
"01010110100000100010011",
"01010110100110100001000",
"01010110101100011111100",
"01010110110010011101111",
"01010110111000011100010",
"01010110111110011010100",
"01010111000100011000101",
"01010111001010010110101",
"01010111010000010100100",
"01010111010110010010010",
"01010111011100010000000",
"01010111100010001101100",
"01010111101000001011000",
"01010111101110001000011",
"01010111110100000101110",
"01010111111010000010111",
"01011000000000000000000",
"01011000000101111100111",
"01011000001011111001110",
"01011000010001110110101",
"01011000010111110011010",
"01011000011101101111110",
"01011000100011101100010",
"01011000101001101000101",
"01011000101111100100111",
"01011000110101100001000",
"01011000111011011101000",
"01011001000001011001000",
"01011001000111010100111",
"01011001001101010000101",
"01011001010011001100010",
"01011001011001000111110",
"01011001011111000011010",
"01011001100100111110100",
"01011001101010111001110",
"01011001110000110100111",
"01011001110110101111111",
"01011001111100101010111",
"01011010000010100101101",
"01011010001000100000011",
"01011010001110011011000",
"01011010010100010101100",
"01011010011010010000000",
"01011010100000001010010",
"01011010100110000100100",
"01011010101011111110101",
"01011010110001111000101",
"01011010110111110010101",
"01011010111101101100011",
"01011011000011100110001",
"01011011001001011111110",
"01011011001111011001010",
"01011011010101010010101",
"01011011011011001100000",
"01011011100001000101010",
"01011011100110111110011",
"01011011101100110111011",
"01011011110010110000010",
"01011011111000101001001",
"01011011111110100001110",
"01011100000100011010011",
"01011100001010010010111",
"01011100010000001011011",
"01011100010110000011101",
"01011100011011111011111",
"01011100100001110100000",
"01011100100111101100000",
"01011100101101100100000",
"01011100110011011011110",
"01011100111001010011100",
"01011100111111001011001",
"01011101000101000010101",
"01011101001010111010001",
"01011101010000110001011",
"01011101010110101000101",
"01011101011100011111110",
"01011101100010010110111",
"01011101101000001101110",
"01011101101110000100101",
"01011101110011111011011",
"01011101111001110010000",
"01011101111111101000100",
"01011110000101011111000",
"01011110001011010101011",
"01011110010001001011101",
"01011110010111000001110",
"01011110011100110111111",
"01011110100010101101110",
"01011110101000100011101",
"01011110101110011001011",
"01011110110100001111001",
"01011110111010000100101",
"01011110111111111010001",
"01011111000101101111100",
"01011111001011100100110",
"01011111010001011010000",
"01011111010111001111000",
"01011111011101000100000",
"01011111100010111001000",
"01011111101000101101110",
"01011111101110100010011",
"01011111110100010111000",
"01011111111010001011100",
"01100000000000000000000",
"01100000000101110100010",
"01100000001011101000100",
"01100000010001011100101",
"01100000010111010000101",
"01100000011101000100101",
"01100000100010111000011",
"01100000101000101100001",
"01100000101110011111110",
"01100000110100010011011",
"01100000111010000110110",
"01100000111111111010001",
"01100001000101101101011",
"01100001001011100000101",
"01100001010001010011101",
"01100001010111000110101",
"01100001011100111001100",
"01100001100010101100010",
"01100001101000011111000",
"01100001101110010001101",
"01100001110100000100001",
"01100001111001110110100",
"01100001111111101000111",
"01100010000101011011000",
"01100010001011001101001",
"01100010010000111111010",
"01100010010110110001001",
"01100010011100100011000",
"01100010100010010100110",
"01100010101000000110011",
"01100010101101110111111",
"01100010110011101001011",
"01100010111001011010110",
"01100010111111001100000",
"01100011000100111101010",
"01100011001010101110010",
"01100011010000011111010",
"01100011010110010000010",
"01100011011100000001000",
"01100011100001110001110",
"01100011100111100010011",
"01100011101101010010111",
"01100011110011000011011",
"01100011111000110011101",
"01100011111110100011111",
"01100100000100010100001",
"01100100001010000100001",
"01100100001111110100001",
"01100100010101100100000",
"01100100011011010011110",
"01100100100001000011100",
"01100100100110110011000",
"01100100101100100010101",
"01100100110010010010000",
"01100100111000000001010",
"01100100111101110000100",
"01100101000011011111101",
"01100101001001001110110",
"01100101001110111101101",
"01100101010100101100100",
"01100101011010011011010",
"01100101100000001010000",
"01100101100101111000101",
"01100101101011100111001",
"01100101110001010101100",
"01100101110111000011110",
"01100101111100110010000",
"01100110000010100000001",
"01100110001000001110001",
"01100110001101111100001",
"01100110010011101010000",
"01100110011001010111110",
"01100110011111000101011",
"01100110100100110011000",
"01100110101010100000100",
"01100110110000001101111",
"01100110110101111011001",
"01100110111011101000011",
"01100111000001010101100",
"01100111000111000010101",
"01100111001100101111100",
"01100111010010011100011",
"01100111011000001001001",
"01100111011101110101110",
"01100111100011100010011",
"01100111101001001110111",
"01100111101110111011010",
"01100111110100100111101",
"01100111111010010011111",
"01101000000000000000000",
"01101000000101101100000",
"01101000001011011000000",
"01101000010001000011111",
"01101000010110101111101",
"01101000011100011011010",
"01101000100010000110111",
"01101000100111110010011",
"01101000101101011101110",
"01101000110011001001001",
"01101000111000110100011",
"01101000111110011111100",
"01101001000100001010101",
"01101001001001110101100",
"01101001001111100000011",
"01101001010101001011010",
"01101001011010110101111",
"01101001100000100000100",
"01101001100110001011000",
"01101001101011110101100",
"01101001110001011111111",
"01101001110111001010001",
"01101001111100110100010",
"01101010000010011110011",
"01101010001101110010010",
"01101010011001000101111",
"01101010100100011001000",
"01101010101111101011111",
"01101010111010111110011",
"01101011000110010000100",
"01101011010001100010010",
"01101011011100110011110",
"01101011101000000100111",
"01101011110011010101101",
"01101011111110100110000",
"01101100001001110110000",
"01101100010101000101110",
"01101100100000010101000",
"01101100101011100100000",
"01101100110110110010110",
"01101101000010000001000",
"01101101001101001111000",
"01101101011000011100101",
"01101101100011101001111",
"01101101101110110110111",
"01101101111010000011011",
"01101110000101001111101",
"01101110010000011011101",
"01101110011011100111001",
"01101110100110110010011",
"01101110110001111101010",
"01101110111101000111111",
"01101111001000010010000",
"01101111010011011011111",
"01101111011110100101011",
"01101111101001101110101",
"01101111110100110111100",
"01110000000000000000000",
"01110000001011001000001",
"01110000010110010000000",
"01110000100001010111100",
"01110000101100011110101",
"01110000110111100101100",
"01110001000010101100000",
"01110001001101110010010",
"01110001011000111000000",
"01110001100011111101100",
"01110001101111000010110",
"01110001111010000111100",
"01110010000101001100000",
"01110010010000010000010",
"01110010011011010100001",
"01110010100110010111101",
"01110010110001011010110",
"01110010111100011101101",
"01110011000111100000001",
"01110011010010100010011",
"01110011011101100100010",
"01110011101000100101110",
"01110011110011100111000",
"01110011111110100111111",
"01110100001001101000100",
"01110100010100101000110",
"01110100011111101000101",
"01110100101010101000010",
"01110100110101100111100",
"01110101000000100110011",
"01110101001011100101000",
"01110101010110100011011",
"01110101100001100001010",
"01110101101100011111000",
"01110101110111011100010",
"01110110000010011001010",
"01110110001101010110000",
"01110110011000010010011",
"01110110100011001110011",
"01110110101110001010001",
"01110110111001000101100",
"01110111000100000000101",
"01110111001110111011011",
"01110111011001110101111",
"01110111100100110000000",
"01110111101111101001111",
"01110111111010100011011",
"01111000000101011100100",
"01111000010000010101011",
"01111000011011001110000",
"01111000100110000110010",
"01111000110000111110001",
"01111000111011110101110",
"01111001000110101101001",
"01111001010001100100001",
"01111001011100011010110",
"01111001100111010001001",
"01111001110010000111001",
"01111001111100111100111",
"01111010000111110010011",
"01111010010010100111100",
"01111010011101011100010",
"01111010101000010000110",
"01111010110011000101000",
"01111010111101111000111",
"01111011001000101100100",
"01111011010011011111110",
"01111011011110010010110",
"01111011101001000101011",
"01111011110011110111110",
"01111011111110101001110",
"01111100001001011011100",
"01111100010100001100111",
"01111100011110111110000",
"01111100101001101110111",
"01111100110100011111011",
"01111100111111001111101",
"01111101001001111111100",
"01111101010100101111001",
"01111101011111011110011",
"01111101101010001101011",
"01111101110100111100001",
"01111101111111101010100",
"01111110001010011000101",
"01111110010101000110011",
"01111110011111110011111",
"01111110101010100001001",
"01111110110101001110000",
"01111110111111111010101",
"01111111001010100110111",
"01111111010101010011000",
"01111111011111111110101",
"01111111101010101010000",
"01111111110101010101001",
"10000000000000000000000",
"10000000001010101010100",
"10000000010101010100110",
"10000000011111111110101",
"10000000101010101000010",
"10000000110101010001101",
"10000000111111111010101",
"10000001001010100011011",
"10000001010101001011111",
"10000001011111110100000",
"10000001101010011011111",
"10000001110101000011100",
"10000001111111101010110",
"10000010001010010001110",
"10000010010100111000100",
"10000010011111011110111",
"10000010101010000101000",
"10000010110100101010110",
"10000010111111010000011",
"10000011001001110101101",
"10000011010100011010100",
"10000011011110111111010",
"10000011101001100011101",
"10000011110100000111110",
"10000011111110101011100",
"10000100001001001111000",
"10000100010011110010010",
"10000100011110010101010",
"10000100101000110111111",
"10000100110011011010010",
"10000100111101111100011",
"10000101001000011110001",
"10000101010010111111101",
"10000101011101100000111",
"10000101101000000001111",
"10000101110010100010100",
"10000101111101000010111",
"10000110000111100011000",
"10000110010010000010111",
"10000110011100100010011",
"10000110100111000001101",
"10000110110001100000101",
"10000110111011111111010",
"10000111000110011101110",
"10000111010000111011111",
"10000111011011011001110",
"10000111100101110111010",
"10000111110000010100101",
"10000111111010110001101",
"10001000000101001110010",
"10001000001111101010110",
"10001000011010000111000",
"10001000100100100010111",
"10001000101110111110100",
"10001000111001011001111",
"10001001000011110100111",
"10001001001110001111101",
"10001001011000101010010",
"10001001100011000100100",
"10001001101101011110011",
"10001001110111111000001",
"10001010000010010001100",
"10001010001100101010101",
"10001010010111000011100",
"10001010100001011100001",
"10001010101011110100100",
"10001010110110001100100",
"10001011000000100100010",
"10001011001010111011110",
"10001011010101010011000",
"10001011011111101010000",
"10001011101010000000101",
"10001011110100010111001",
"10001011111110101101010",
"10001100001001000011001",
"10001100010011011000110",
"10001100011101101110000",
"10001100101000000011001",
"10001100110010010111111",
"10001100111100101100100",
"10001101000111000000110",
"10001101010001010100110",
"10001101011011101000100",
"10001101100101111011111",
"10001101110000001111001",
"10001101111010100010000",
"10001110000100110100110",
"10001110001111000111001",
"10001110011001011001010",
"10001110100011101011001",
"10001110101101111100101",
"10001110111000001110000",
"10001111000010011111001",
"10001111001100101111111",
"10001111010111000000011",
"10001111100001010000110",
"10001111101011100000110",
"10001111110101110000100",
"10010000000000000000000",
"10010000001010001111010",
"10010000010100011110001",
"10010000011110101100111",
"10010000101000111011011",
"10010000110011001001100",
"10010000111101010111011",
"10010001000111100101001",
"10010001010001110010100",
"10010001011011111111101",
"10010001100110001100100",
"10010001110000011001001",
"10010001111010100101100",
"10010010000100110001101",
"10010010001110111101100",
"10010010011001001001000",
"10010010100011010100011",
"10010010101101011111100",
"10010010110111101010010",
"10010011000001110100111",
"10010011001011111111001",
"10010011010110001001010",
"10010011100000010011000",
"10010011101010011100100",
"10010011110100100101111",
"10010011111110101110111",
"10010100001000110111101",
"10010100010011000000001",
"10010100011101001000011",
"10010100100111010000100",
"10010100110001011000010",
"10010100111011011111110",
"10010101000101100111000",
"10010101001111101110000",
"10010101011001110100110",
"10010101100011111011010",
"10010101101110000001100",
"10010101111000000111100",
"10010110000010001101010",
"10010110001100010010110",
"10010110010110011000000",
"10010110100000011101000",
"10010110101010100001110",
"10010110110100100110001",
"10010110111110101010011",
"10010111001000101110011",
"10010111010010110010001",
"10010111011100110101101",
"10010111100110111000111",
"10010111110000111011111",
"10010111111010111110110",
"10011000000101000001010",
"10011000001111000011100",
"10011000011001000101100",
"10011000100011000111010",
"10011000101101001000110",
"10011000110111001010000",
"10011001000001001011001",
"10011001001011001011111",
"10011001010101001100011",
"10011001011111001100110",
"10011001101001001100110",
"10011001110011001100101",
"10011001111101001100001",
"10011010000111001011100",
"10011010010001001010100",
"10011010011011001001011",
"10011010100101001000000",
"10011010101111000110011",
"10011010111001000100011",
"10011011000011000010010",
"10011011001100111111111",
"10011011010110111101010",
"10011011100000111010100",
"10011011101010110111011",
"10011011110100110100000",
"10011011111110110000100",
"10011100001000101100101",
"10011100010010101000101",
"10011100011100100100010",
"10011100100110011111110",
"10011100110000011011000",
"10011100111010010110000",
"10011101000100010000110",
"10011101001110001011010",
"10011101011000000101100",
"10011101100001111111100",
"10011101101011111001010",
"10011101110101110010111",
"10011101111111101100010",
"10011110001001100101010",
"10011110010011011110001",
"10011110011101010110110",
"10011110100111001111001",
"10011110110001000111010",
"10011110111010111111001",
"10011111000100110110111",
"10011111001110101110010",
"10011111011000100101100",
"10011111100010011100100",
"10011111101100010011010",
"10011111110110001001110",
"10100000000000000000000",
"10100000001001110110000",
"10100000010011101011111",
"10100000011101100001011",
"10100000100111010110110",
"10100000110001001011111",
"10100000111011000000110",
"10100001000100110101011",
"10100001001110101001110",
"10100001011000011110000",
"10100001100010010001111",
"10100001101100000101101",
"10100001110101111001001",
"10100001111111101100011",
"10100010001001011111011",
"10100010010011010010010",
"10100010011101000100110",
"10100010100110110111001",
"10100010110000101001010",
"10100010111010011011001",
"10100011000100001100110",
"10100011001101111110010",
"10100011010111101111011",
"10100011100001100000011",
"10100011101011010001001",
"10100011110101000001101",
"10100011111110110010000",
"10100100001000100010000",
"10100100010010010001111",
"10100100011100000001100",
"10100100100101110000111",
"10100100101111100000000",
"10100100111001001111000",
"10100101000010111101101",
"10100101001100101100001",
"10100101010110011010100",
"10100101100000001000100",
"10100101101001110110010",
"10100101110011100011111",
"10100101111101010001010",
"10100110000110111110011",
"10100110010000101011011",
"10100110011010011000000",
"10100110100100000100100",
"10100110101101110000110",
"10100110110111011100110",
"10100111000001001000101",
"10100111001010110100001",
"10100111010100011111100",
"10100111011110001010110",
"10100111100111110101101",
"10100111110001100000011",
"10100111111011001010111",
"10101000000100110101001",
"10101000001110011111001",
"10101000011000001001000",
"10101000100001110010100",
"10101000101011011100000",
"10101000110101000101001",
"10101000111110101110000",
"10101001001000010110110",
"10101001010001111111010",
"10101001011011100111101",
"10101001100101001111101",
"10101001101110110111100",
"10101001111000011111001",
"10101010000010000110101",
"10101010001011101101110",
"10101010010101010100110",
"10101010011110111011100",
"10101010101000100010001",
"10101010110010001000100",
"10101010111011101110101",
"10101011000101010100100",
"10101011001110111010001",
"10101011011000011111101",
"10101011100010000100111",
"10101011101011101010000",
"10101011110101001110110",
"10101011111110110011011",
"10101100001000010111111",
"10101100010001111100000",
"10101100011011100000000",
"10101100100101000011110",
"10101100101110100111010",
"10101100111000001010101",
"10101101000001101101110",
"10101101001011010000101",
"10101101010100110011011",
"10101101011110010101111",
"10101101100111111000001",
"10101101110001011010010",
"10101101111010111100001",
"10101110000100011101110",
"10101110001101111111001",
"10101110010111100000011",
"10101110100001000001011",
"10101110101010100010001",
"10101110110100000010110",
"10101110111101100011001",
"10101111000111000011011",
"10101111010000100011010",
"10101111011010000011000",
"10101111100011100010101",
"10101111101101000001111",
"10101111110110100001000",
"10110000000000000000000",
"10110000001001011110101",
"10110000010010111101010",
"10110000011100011011100",
"10110000100101111001101",
"10110000101111010111100",
"10110000111000110101001",
"10110001000010010010101",
"10110001001011101111111",
"10110001010101001100111",
"10110001011110101001110",
"10110001101000000110011",
"10110001110001100010111",
"10110001111010111111000",
"10110010000100011011001",
"10110010001101110110111",
"10110010010111010010100",
"10110010100000101101111",
"10110010101010001001001",
"10110010110011100100001",
"10110010111100111110111",
"10110011000110011001100",
"10110011001111110011111",
"10110011011001001110001",
"10110011100010101000001",
"10110011101100000001111",
"10110011110101011011100",
"10110011111110110100111",
"10110100001000001110000",
"10110100010001100111000",
"10110100011010111111110",
"10110100100100011000010",
"10110100101101110000101",
"10110100110111001000111",
"10110101000000100000110",
"10110101001001111000100",
"10110101010011010000001",
"10110101011100100111100",
"10110101100101111110101",
"10110101101111010101101",
"10110101111000101100011",
"10110110000010000010111",
"10110110001011011001010",
"10110110010100101111011",
"10110110011110000101011",
"10110110100111011011001",
"10110110110000110000110",
"10110110111010000110000",
"10110111000011011011010",
"10110111001100110000010",
"10110111010110000101000",
"10110111011111011001100",
"10110111101000101101111",
"10110111110010000010001",
"10110111111011010110000",
"10111000000100101001111",
"10111000001101111101011",
"10111000010111010000111",
"10111000100000100100000",
"10111000101001110111000",
"10111000110011001001110",
"10111000111100011100011",
"10111001000101101110110",
"10111001001111000001000",
"10111001011000010011000",
"10111001100001100100111",
"10111001101010110110100",
"10111001110100000111111",
"10111001111101011001001",
"10111010000110101010010",
"10111010001111111011000",
"10111010011001001011110",
"10111010100010011100001",
"10111010101011101100100",
"10111010110100111100100",
"10111010111110001100011",
"10111011000111011100001",
"10111011010000101011101",
"10111011011001111010111",
"10111011100011001010000",
"10111011101100011000111",
"10111011110101100111101",
"10111011111110110110001",
"10111100001000000100100",
"10111100010001010010101",
"10111100011010100000101",
"10111100100011101110011",
"10111100101100111100000",
"10111100110110001001011",
"10111100111111010110100",
"10111101001000100011100",
"10111101010001110000011",
"10111101011010111101000",
"10111101100100001001011",
"10111101101101010101101",
"10111101110110100001110",
"10111101111111101101101",
"10111110001000111001010",
"10111110010010000100110",
"10111110011011010000001",
"10111110100100011011001",
"10111110101101100110001",
"10111110110110110000111",
"10111110111111111011011",
"10111111001001000101110",
"10111111010010001111111",
"10111111011011011001111",
"10111111100100100011110",
"10111111101101101101011",
"10111111110110110110110",
"11000000000000000000000",
"11000000001001001001000",
"11000000010010010001111",
"11000000011011011010101",
"11000000100100100011000",
"11000000101101101011011",
"11000000110110110011100",
"11000000111111111011011",
"11000001001001000011001",
"11000001010010001010110",
"11000001011011010010001",
"11000001100100011001010",
"11000001101101100000010",
"11000001110110100111001",
"11000001111111101101110",
"11000010001000110100010",
"11000010010001111010100",
"11000010011011000000101",
"11000010100100000110100",
"11000010101101001100010",
"11000010110110010001110",
"11000010111111010111001",
"11000011001000011100010",
"11000011010001100001010",
"11000011011010100110001",
"11000011100011101010110",
"11000011101100101111001",
"11000011110101110011011",
"11000011111110110111100",
"11000100000111111011011",
"11000100010000111111001",
"11000100011010000010101",
"11000100100011000110000",
"11000100101100001001001",
"11000100110101001100001",
"11000100111110001111000",
"11000101000111010001101",
"11000101010000010100000",
"11000101011001010110010",
"11000101100010011000011",
"11000101101011011010010",
"11000101110100011100000",
"11000101111101011101101",
"11000110000110011111000",
"11000110001111100000001",
"11000110011000100001001",
"11000110100001100010000",
"11000110101010100010101",
"11000110110011100011001",
"11000110111100100011011",
"11000111000101100011100",
"11000111001110100011100",
"11000111010111100011010",
"11000111100000100010111",
"11000111101001100010010",
"11000111110010100001100",
"11000111111011100000100",
"11001000000100011111011",
"11001000001101011110001",
"11001000010110011100101",
"11001000011111011011000",
"11001000101000011001001",
"11001000110001010111001",
"11001000111010010101000",
"11001001000011010010101",
"11001001001100010000000",
"11001001010101001101011",
"11001001011110001010100",
"11001001100111000111011",
"11001001110000000100001",
"11001001111001000000110",
"11001010000001111101001",
"11001010001010111001011",
"11001010010011110101100",
"11001010011100110001011",
"11001010100101101101001",
"11001010101110101000101",
"11001010110111100100000",
"11001011000000011111010",
"11001011001001011010010",
"11001011010010010101001",
"11001011011011001111110",
"11001011100100001010010",
"11001011101101000100101",
"11001011110101111110110",
"11001011111110111000110",
"11001100000111110010100",
"11001100010000101100010",
"11001100011001100101101",
"11001100100010011111000",
"11001100101011011000001",
"11001100110100010001000",
"11001100111101001001111",
"11001101000110000010011",
"11001101001110111010111",
"11001101010111110011001",
"11001101100000101011010",
"11001101101001100011001",
"11001101110010011010111",
"11001101111011010010100",
"11001110000100001001111",
"11001110001101000001001",
"11001110010101111000010",
"11001110011110101111001",
"11001110100111100101111",
"11001110110000011100100",
"11001110111001010010111",
"11001111000010001001001",
"11001111001010111111001",
"11001111010011110101000",
"11001111011100101010110",
"11001111100101100000011",
"11001111101110010101110",
"11001111110111001010111",
"11010000000000000000000",
"11010000001000110100111",
"11010000010001101001101",
"11010000011010011110001",
"11010000100011010010100",
"11010000101100000110110",
"11010000110100111010110",
"11010000111101101110101",
"11010001000110100010011",
"11010001001111010101111",
"11010001011000001001010",
"11010001100000111100100",
"11010001101001101111100",
"11010001110010100010011",
"11010001111011010101001",
"11010010000100000111101",
"11010010001100111010000",
"11010010010101101100010",
"11010010011110011110010",
"11010010100111010000001",
"11010010110000000001111",
"11010010111000110011100",
"11010011000001100100111",
"11010011001010010110000",
"11010011010011000111001",
"11010011011011111000000",
"11010011100100101000110",
"11010011101101011001010",
"11010011110110001001110",
"11010011111110111010000",
"11010100000111101010000",
"11010100010000011010000",
"11010100011001001001110",
"11010100100001111001010",
"11010100101010101000110",
"11010100110011011000000",
"11010100111100000111000",
"11010101000100110110000",
"11010101001101100100110",
"11010101010110010011011",
"11010101011111000001110",
"11010101100111110000001",
"11010101110000011110010",
"11010101111001001100001",
"11010110000001111010000",
"11010110001010100111101",
"11010110010011010101001",
"11010110011100000010011",
"11010110100100101111100",
"11010110101101011100100",
"11010110110110001001011",
"11010110111110110110000",
"11010111000111100010100",
"11010111010000001110111",
"11010111011000111011001",
"11010111100001100111001",
"11010111101010010011000",
"11010111110010111110110",
"11010111111011101010010",
"11011000000100010101101",
"11011000001101000000111",
"11011000010101101100000",
"11011000011110010110111",
"11011000100111000001101",
"11011000101111101100010",
"11011000111000010110101",
"11011001000001000000111",
"11011001001001101011000",
"11011001010010010101000",
"11011001011010111110110",
"11011001100011101000100",
"11011001101100010001111",
"11011001110100111011010",
"11011001111101100100011",
"11011010000110001101011",
"11011010001110110110010",
"11011010010111011111000",
"11011010100000000111100",
"11011010101000101111111",
"11011010110001011000001",
"11011010111010000000010",
"11011011000010101000001",
"11011011001011001111111",
"11011011010011110111100",
"11011011011100011110111",
"11011011100101000110010",
"11011011101101101101011",
"11011011110110010100010",
"11011011111110111011001",
"11011100000111100001110",
"11011100010000001000010",
"11011100011000101110101",
"11011100100001010100111",
"11011100101001111010111",
"11011100110010100000110",
"11011100111011000110100",
"11011101000011101100001",
"11011101001100010001100",
"11011101010100110110110",
"11011101011101011011111",
"11011101100110000000111",
"11011101101110100101101",
"11011101110111001010011",
"11011101111111101110111",
"11011110001000010011001",
"11011110010000110111011",
"11011110011001011011011",
"11011110100001111111010",
"11011110101010100011000",
"11011110110011000110101",
"11011110111011101010000",
"11011111000100001101011",
"11011111001100110000011",
"11011111010101010011011",
"11011111011101110110010",
"11011111100110011000111",
"11011111101110111011011",
"11011111110111011101110",
"11100000000000000000000",
"11100000001000100010000",
"11100000010001000011111",
"11100000011001100101110",
"11100000100010000111010",
"11100000101010101000110",
"11100000110011001010000",
"11100000111011101011010",
"11100001000100001100010",
"11100001001100101101000",
"11100001010101001101110",
"11100001011101101110010",
"11100001100110001110101",
"11100001101110101110111",
"11100001110111001111000",
"11100001111111101111000",
"11100010001000001110110",
"11100010010000101110011",
"11100010011001001101111",
"11100010100001101101010",
"11100010101010001100100",
"11100010110010101011100",
"11100010111011001010011",
"11100011000011101001001",
"11100011001100000111110",
"11100011010100100110010",
"11100011011101000100100",
"11100011100101100010101",
"11100011101110000000110",
"11100011110110011110100",
"11100011111110111100010",
"11100100000111011001111",
"11100100001111110111010",
"11100100011000010100100",
"11100100100000110001101",
"11100100101001001110101",
"11100100110001101011011",
"11100100111010001000001",
"11100101000010100100101",
"11100101001011000001000",
"11100101010011011101010",
"11100101011011111001011",
"11100101100100010101010",
"11100101101100110001001",
"11100101110101001100110",
"11100101111101101000010",
"11100110000110000011101",
"11100110001110011110111",
"11100110010110111001111",
"11100110011111010100111",
"11100110100111101111101",
"11100110110000001010010",
"11100110111000100100110",
"11100111000000111111000",
"11100111001001011001010",
"11100111010001110011010",
"11100111011010001101010",
"11100111100010100111000",
"11100111101011000000101",
"11100111110011011010000",
"11100111111011110011011",
"11101000000100001100100",
"11101000001100100101101",
"11101000010100111110100",
"11101000011101010111010",
"11101000100101101111111",
"11101000101110001000010",
"11101000110110100000101",
"11101000111110111000110",
"11101001000111010000110",
"11101001001111101000101",
"11101001011000000000011",
"11101001100000011000000",
"11101001101000101111100",
"11101001110001000110110",
"11101001111001011110000",
"11101010000001110101000",
"11101010001010001011111",
"11101010010010100010101",
"11101010011010111001010",
"11101010100011001111101",
"11101010101011100110000",
"11101010110011111100001",
"11101010111100010010010",
"11101011000100101000001",
"11101011001100111101111",
"11101011010101010011100",
"11101011011101101000111",
"11101011100101111110010",
"11101011101110010011011",
"11101011110110101000100",
"11101011111110111101011",
"11101100000111010010001",
"11101100001111100110110",
"11101100010111111011010",
"11101100100000001111101",
"11101100101000100011110",
"11101100110000110111111",
"11101100111001001011110",
"11101101000001011111100",
"11101101001001110011001",
"11101101010010000110101",
"11101101011010011010000",
"11101101100010101101010",
"11101101101011000000010",
"11101101110011010011010",
"11101101111011100110000",
"11101110000011111000110",
"11101110001100001011010",
"11101110010100011101101",
"11101110011100101111111",
"11101110100101000010000",
"11101110101101010011111",
"11101110110101100101110",
"11101110111101110111011",
"11101111000110001001000",
"11101111001110011010011",
"11101111010110101011101",
"11101111011110111100110",
"11101111100111001101110",
"11101111101111011110101",
"11101111110111101111011",
"11110000000000000000000",
"11110000001000010000011",
"11110000010000100000110",
"11110000011000110000111",
"11110000100001000000111",
"11110000101001010000111",
"11110000110001100000101",
"11110000111001110000010",
"11110001000001111111110",
"11110001001010001111000",
"11110001010010011110010",
"11110001011010101101011",
"11110001100010111100010",
"11110001101011001011001",
"11110001110011011001110",
"11110001111011101000010",
"11110010000011110110110",
"11110010001100000101000",
"11110010010100010011001",
"11110010011100100001001",
"11110010100100101110111",
"11110010101100111100101",
"11110010110101001010010",
"11110010111101010111110",
"11110011000101100101000",
"11110011001101110010001",
"11110011010101111111010",
"11110011011110001100001",
"11110011100110011000111",
"11110011101110100101100",
"11110011110110110010000",
"11110011111110111110011",
"11110100000111001010101",
"11110100001111010110110",
"11110100010111100010110",
"11110100011111101110101",
"11110100100111111010010",
"11110100110000000101111",
"11110100111000010001010",
"11110101000000011100101",
"11110101001000100111110",
"11110101010000110010110",
"11110101011000111101101",
"11110101100001001000100",
"11110101101001010011001",
"11110101110001011101101",
"11110101111001101000000",
"11110110000001110010010",
"11110110001001111100010",
"11110110010010000110010",
"11110110011010010000001",
"11110110100010011001111",
"11110110101010100011011",
"11110110110010101100111",
"11110110111010110110001",
"11110111000010111111011",
"11110111001011001000011",
"11110111010011010001010",
"11110111011011011010001",
"11110111100011100010110",
"11110111101011101011010",
"11110111110011110011101",
"11110111111011111011111",
"11111000000100000100000",
"11111000001100001100000",
"11111000010100010011111",
"11111000011100011011101",
"11111000100100100011010",
"11111000101100101010110",
"11111000110100110010000",
"11111000111100111001010",
"11111001000101000000011",
"11111001001101000111010",
"11111001010101001110001",
"11111001011101010100110",
"11111001100101011011011",
"11111001101101100001110",
"11111001110101101000001",
"11111001111101101110010",
"11111010000101110100010",
"11111010001101111010010",
"11111010010110000000000",
"11111010011110000101101",
"11111010100110001011001",
"11111010101110010000101",
"11111010110110010101111",
"11111010111110011011000",
"11111011000110100000000",
"11111011001110100100111",
"11111011010110101001101",
"11111011011110101110010",
"11111011100110110010110",
"11111011101110110111001",
"11111011110110111011011",
"11111011111110111111100",
"11111100000111000011100",
"11111100001111000111010",
"11111100010111001011000",
"11111100011111001110101",
"11111100100111010010001",
"11111100101111010101100",
"11111100110111011000101",
"11111100111111011011110",
"11111101000111011110110",
"11111101001111100001100",
"11111101010111100100010",
"11111101011111100110111",
"11111101100111101001010",
"11111101101111101011101",
"11111101110111101101111",
"11111101111111101111111",
"11111110000111110001111",
"11111110001111110011101",
"11111110010111110101011",
"11111110011111110111000",
"11111110100111111000011",
"11111110101111111001110",
"11111110110111111010111",
"11111110111111111100000",
"11111111000111111100111",
"11111111001111111101110",
"11111111010111111110011",
"11111111011111111111000",
"11111111100111111111011",
"11111111101111111111110",
"11111111110111111111111");
  constant rom2 : rom_t :=("00000000000000000000000",
"11111111110000000000110",
"11111111100000000011000",
"11111111010000000110110",
"11111111000000001100000",
"11111110110000010010110",
"11111110100000011011000",
"11111110010000100100101",
"11111110000000101111111",
"11111101110000111100100",
"11111101100001001010101",
"11111101010001011010001",
"11111101000001101011000",
"11111100110001111101100",
"11111100100010010001100",
"11111100010010100110111",
"11111100000010111101101",
"11111011110011010110000",
"11111011100011101111100",
"11111011010100001010110",
"11111011000100100111010",
"11111010110101000101011",
"11111010100101100100110",
"11111010010110000101100",
"11111010000110101000000",
"11111001110111001011101",
"11111001100111110000101",
"11111001011000010111001",
"11111001001000111111001",
"11111000111001101000100",
"11111000101010010011000",
"11111000011010111111001",
"11111000001011101100110",
"11110111111100011011100",
"11110111101101001011110",
"11110111011101111101100",
"11110111001110110000100",
"11110110111111100100111",
"11110110110000011010101",
"11110110100001010001111",
"11110110010010001010011",
"11110110000011000100001",
"11110101110011111111100",
"11110101100100111100000",
"11110101010101111010001",
"11110101000110111001011",
"11110100110111111010000",
"11110100101000111100000",
"11110100011001111111011",
"11110100001011000011111",
"11110011111100001010000",
"11110011101101010001001",
"11110011011110011010000",
"11110011001111100100000",
"11110011000000101111010",
"11110010110001111100000",
"11110010100011001001110",
"11110010010100011001001",
"11110010000101101001101",
"11110001110110111011011",
"11110001101000001110101",
"11110001011001100011001",
"11110001001010111001000",
"11110000111100010000001",
"11110000101101101000011",
"11110000011111000010000",
"11110000010000011100111",
"11110000000001111001010",
"11101111110011010110110",
"11101111100100110101100",
"11101111010110010101101",
"11101111000111110111000",
"11101110111001011001101",
"11101110101010111101010",
"11101110011100100010100",
"11101110001110001000110",
"11101101111111110000011",
"11101101110001011001011",
"11101101100011000011100",
"11101101010100101111000",
"11101101000110011011101",
"11101100111000001001100",
"11101100101001111000101",
"11101100011011101000111",
"11101100001101011010101",
"11101011111111001101011",
"11101011110001000001011",
"11101011100010110110110",
"11101011010100101101001",
"11101011000110100101000",
"11101010111000011110000",
"11101010101010011000001",
"11101010011100010011011",
"11101010001110001111111",
"11101010000000001101111",
"11101001110010001100101",
"11101001100100001101000",
"11101001010110001110010",
"11101001001000010000111",
"11101000111010010100101",
"11101000101100011001110",
"11101000011110011111111",
"11101000010000100111001",
"11101000000010101111110",
"11100111110100111001100",
"11100111100111000100011",
"11100111011001010000100",
"11100111001011011101110",
"11100110111101101100001",
"11100110101111111011101",
"11100110100010001100011",
"11100110010100011110011",
"11100110000110110001011",
"11100101111001000101101",
"11100101101011011011000",
"11100101011101110001100",
"11100101010000001001001",
"11100101000010100010000",
"11100100110100111011110",
"11100100100111010111001",
"11100100011001110011011",
"11100100001100010000101",
"11100011111110101111010",
"11100011110001001110111",
"11100011100011101111100",
"11100011010110010001101",
"11100011001000110100101",
"11100010111011011000101",
"11100010101101111110000",
"11100010100000100100011",
"11100010010011001100000",
"11100010000101110100100",
"11100001111000011110001",
"11100001101011001001000",
"11100001011101110100111",
"11100001010000100010001",
"11100001000011010000001",
"11100000110101111111100",
"11100000101000101111111",
"11100000011011100001011",
"11100000001110010011110",
"11100000000001000111011",
"11011111110011111100001",
"11011111100110110001111",
"11011111011001101000110",
"11011111001100100000110",
"11011110111111011001110",
"11011110110010010011111",
"11011110100101001110111",
"11011110011000001011001",
"11011110001011001000100",
"11011101111110000111000",
"11011101110001000110011",
"11011101100100000110110",
"11011101010111001000100",
"11011101001010001011001",
"11011100111101001110101",
"11011100110000010011011",
"11011100100011011001001",
"11011100010110011111111",
"11011100001001100111110",
"11011011111100110000110",
"11011011101111111010101",
"11011011100011000101110",
"11011011010110010001101",
"11011011001001011110111",
"11011010111100101100111",
"11011010101111111100000",
"11011010100011001100001",
"11011010010110011101100",
"11011010001001101111101",
"11011001111101000010110",
"11011001110000010111000",
"11011001100011101100010",
"11011001010111000010100",
"11011001001010011001110",
"11011000111101110010010",
"11011000110001001011100",
"11011000100100100101101",
"11011000011000000001001",
"11011000001011011101011",
"11010111111110111010110",
"11010111110010011001001",
"11010111100101111000011",
"11010111011001011000101",
"11010111001100111010000",
"11010111000000011100010",
"11010110110011111111101",
"11010110100111100011111",
"11010110011011001001001",
"11010110001110101111010",
"11010110000010010110100",
"11010101110101111110111",
"11010101101001101000000",
"11010101011101010010000",
"11010101010000111101001",
"11010101000100101001010",
"11010100111000010110011",
"11010100101100000100011",
"11010100011111110011011",
"11010100010011100011011",
"11010100000111010100001",
"11010011111011000110001",
"11010011101110111000110",
"11010011100010101100101",
"11010011010110100001100",
"11010011001010010111001",
"11010010111110001101110",
"11010010110010000101010",
"11010010100101111101111",
"11010010011001110111011",
"11010010001101110001101",
"11010010000001101101000",
"11010001110101101001011",
"11010001101001100110101",
"11010001011101100100101",
"11010001010001100011101",
"11010001000101100011110",
"11010000111001100100110",
"11010000101101100110101",
"11010000100001101001100",
"11010000010101101101000",
"11010000001001110001101",
"11001111111101110111011",
"11001111110001111101110",
"11001111100110000101001",
"11001111011010001101011",
"11001111001110010110101",
"11001111000010100000110",
"11001110110110101011110",
"11001110101010110111101",
"11001110011111000100100",
"11001110010011010010010",
"11001110000111100001000",
"11001101111011110000011",
"11001101110000000000111",
"11001101100100010010001",
"11001101011000100100100",
"11001101001100110111100",
"11001101000001001011011",
"11001100110101100000011",
"11001100101001110110001",
"11001100011110001100110",
"11001100010010100100010",
"11001100000110111100110",
"11001011111011010110001",
"11001011101111110000010",
"11001011100100001011011",
"11001011011000100111010",
"11001011001101000100001",
"11001011000001100001110",
"11001010110110000000001",
"11001010101010011111101",
"11001010011111000000000",
"11001010010011100001000",
"11001010001000000011001",
"11001001111100100101110",
"11001001110001001001101",
"11001001100101101110001",
"11001001011010010011101",
"11001001001110111010000",
"11001001000011100000111",
"11001000111000001001000",
"11001000101100110001110",
"11001000100001011011011",
"11001000010110000110000",
"11001000001010110001011",
"11000111111111011101100",
"11000111110100001010101",
"11000111101000111000100",
"11000111011101100111010",
"11000111010010010110111",
"11000111000111000111001",
"11000110111011111000011",
"11000110110000101010100",
"11000110100101011101011",
"11000110011010010001001",
"11000110001111000101101",
"11000110000011111011000",
"11000101111000110001001",
"11000101101101101000010",
"11000101100010100000000",
"11000101010111011000101",
"11000101001100010010001",
"11000101000001001100011",
"11000100110110000111100",
"11000100101011000011100",
"11000100100000000000001",
"11000100010100111101110",
"11000100001001111100000",
"11000011111110111011001",
"11000011110011111011000",
"11000011101000111011110",
"11000011011101111101011",
"11000011010010111111110",
"11000011001000000010111",
"11000010111101000110111",
"11000010110010001011100",
"11000010100111010001000",
"11000010011100010111011",
"11000010010001011110100",
"11000010000110100110100",
"11000001111011101111001",
"11000001110000111000101",
"11000001100110000010110",
"11000001011011001101110",
"11000001010000011001101",
"11000001000101100110010",
"11000000111010110011101",
"11000000110000000001110",
"11000000100101010000110",
"11000000011010100000011",
"11000000001111110000111",
"11000000000101000010001",
"10111111111010010100001",
"10111111101111100111001",
"10111111100100111010100",
"10111111011010001110111",
"10111111001111100100000",
"10111111000100111001110",
"10111110111010010000011",
"10111110101111100111111",
"10111110100101000000000",
"10111110011010011000111",
"10111110001111110010100",
"10111110000101001101000",
"10111101111010101000001",
"10111101110000000011111",
"10111101100101100000101",
"10111101011010111110000",
"10111101010000011100001",
"10111101000101111011001",
"10111100111011011010101",
"10111100110000111011001",
"10111100100110011100001",
"10111100011011111110000",
"10111100010001100000101",
"10111100000111000100001",
"10111011111100101000000",
"10111011110010001101000",
"10111011100111110010100",
"10111011011101011000111",
"10111011010010111111111",
"10111011001000100111100",
"10111010111110001111111",
"10111010110011111001001",
"10111010101001100011000",
"10111010011111001101110",
"10111010010100111001010",
"10111010001010100101010",
"10111010000000010010000",
"10111001110101111111101",
"10111001101011101101110",
"10111001100001011100111",
"10111001010111001100100",
"10111001001100111100111",
"10111001000010101110000",
"10111000111000011111110",
"10111000101110010010011",
"10111000100100000101101",
"10111000011001111001101",
"10111000001111101110001",
"10111000000101100011101",
"10110111111011011001101",
"10110111110001010000011",
"10110111100111000111110",
"10110111011101000000000",
"10110111010010111000111",
"10110111001000110010011",
"10110110111110101100110",
"10110110110100100111110",
"10110110101010100011011",
"10110110100000011111101",
"10110110010110011100110",
"10110110001100011010100",
"10110110000010011000111",
"10110101111000011000000",
"10110101101110010111110",
"10110101100100011000001",
"10110101011010011001010",
"10110101010000011011010",
"10110101000110011101101",
"10110100111100100000111",
"10110100110010100100110",
"10110100101000101001010",
"10110100011110101110100",
"10110100010100110100100",
"10110100001010111011001",
"10110100000001000010010",
"10110011110111001010011",
"10110011101101010010110",
"10110011100011011100000",
"10110011011001100110000",
"10110011001111110000101",
"10110011000101111011111",
"10110010111100000111110",
"10110010110010010100011",
"10110010101000100001110",
"10110010011110101111100",
"10110010010100111110001",
"10110010001011001101011",
"10110010000001011101010",
"10110001110111101101111",
"10110001101101111111000",
"10110001100100010000111",
"10110001011010100011011",
"10110001010000110110110",
"10110001000111001010100",
"10110000111101011111000",
"10110000110011110100001",
"10110000101010001001111",
"10110000100000100000010",
"10110000010110110111011",
"10110000001101001110111",
"10110000000011100111010",
"10101111111010000000011",
"10101111110000011010000",
"10101111100110110100001",
"10101111011101001111001",
"10101111010011101010101",
"10101111001010000110110",
"10101111000000100011110",
"10101110110111000001001",
"10101110101101011111010",
"10101110100011111101111",
"10101110011010011101010",
"10101110010000111101001",
"10101110000111011101111",
"10101101111101111111000",
"10101101110100100000111",
"10101101101011000011011",
"10101101100001100110011",
"10101101011000001010010",
"10101101001110101110100",
"10101101000101010011100",
"10101100111011111001001",
"10101100110010011111011",
"10101100101001000110001",
"10101100011111101101101",
"10101100010110010101101",
"10101100001100111110010",
"10101100000011100111101",
"10101011111010010001100",
"10101011110000111100001",
"10101011100111100111001",
"10101011011110010011000",
"10101011010100111111011",
"10101011001011101100010",
"10101011000010011001111",
"10101010111001001000000",
"10101010101111110110101",
"10101010100110100110001",
"10101010011101010110001",
"10101010010100000110110",
"10101010001010110111111",
"10101010000001101001101",
"10101001111000011011111",
"10101001101111001111000",
"10101001100110000010011",
"10101001011100110110101",
"10101001010011101011011",
"10101001001010100000110",
"10101001000001010110110",
"10101000111000001101010",
"10101000101111000100011",
"10101000100101111100000",
"10101000011100110100011",
"10101000010011101101010",
"10101000001010100110110",
"10101000000001100000110",
"10100111111000011011100",
"10100111101111010110101",
"10100111100110010010100",
"10100111011101001110111",
"10100111010100001011111",
"10100111001011001001011",
"10100111000010000111100",
"10100110111001000110010",
"10100110110000000101101",
"10100110100111000101011",
"10100110011110000101111",
"10100110010101000110111",
"10100110001100001000100",
"10100110000011001010101",
"10100101111010001101010",
"10100101110001010000100",
"10100101101000010100011",
"10100101011111011000111",
"10100101010110011101111",
"10100101001101100011011",
"10100101000100101001100",
"10100100111011110000010",
"10100100110010110111100",
"10100100101001111111010",
"10100100100001000111110",
"10100100011000010000101",
"10100100001111011010010",
"10100100000110100100001",
"10100011111101101110110",
"10100011110100111010000",
"10100011101100000101110",
"10100011100011010010000",
"10100011011010011110111",
"10100011010001101100010",
"10100011001000111010010",
"10100011000000001000101",
"10100010110111010111110",
"10100010101110100111010",
"10100010100101110111100",
"10100010011101001000010",
"10100010010100011001100",
"10100010001011101011010",
"10100010000010111101101",
"10100001111010010000011",
"10100001110001100011110",
"10100001101000110111110",
"10100001100000001100010",
"10100001010111100001010",
"10100001001110110110111",
"10100001000110001101001",
"10100000111101100011101",
"10100000110100111010111",
"10100000101100010010101",
"10100000100011101010111",
"10100000011011000011101",
"10100000010010011101000",
"10100000001001110111000",
"10100000000001010001011",
"10011111111000101100010",
"10011111110000000111110",
"10011111100111100011101",
"10011111011111000000010",
"10011111010110011101011",
"10011111001101111010111",
"10011111000101011001000",
"10011110111100110111101",
"10011110110100010110111",
"10011110101011110110100",
"10011110100011010110110",
"10011110011010110111011",
"10011110010010011000101",
"10011110001001111010011",
"10011110000001011100110",
"10011101111000111111100",
"10011101110000100010110",
"10011101101000000110101",
"10011101011111101011000",
"10011101010111001111111",
"10011101001110110101011",
"10011101000110011011001",
"10011100111110000001101",
"10011100110101101000100",
"10011100101101010000000",
"10011100100100111000000",
"10011100011100100000010",
"10011100010100001001010",
"10011100001011110010110",
"10011100000011011100110",
"10011011111011000111011",
"10011011110010110010010",
"10011011101010011101110",
"10011011100010001001110",
"10011011011001110110010",
"10011011010001100011011",
"10011011001001010000110",
"10011011000000111110110",
"10011010111000101101011",
"10011010110000011100010",
"10011010101000001011111",
"10011010011111111011110",
"10011010010111101100011",
"10011010001111011101010",
"10011010000111001110111",
"10011001111111000000110",
"10011001110110110011010",
"10011001101110100110010",
"10011001100110011001101",
"10011001011110001101101",
"10011001010110000010001",
"10011001001101110111001",
"10011001000101101100011",
"10011000111101100010011",
"10011000110101011000110",
"10011000101101001111110",
"10011000100101000111001",
"10011000011100111110111",
"10011000010100110111010",
"10011000001100110000000",
"10011000000100101001011",
"10010111111100100011001",
"10010111110100011101100",
"10010111101100011000010",
"10010111100100010011100",
"10010111011100001111010",
"10010111010100001011011",
"10010111001100001000001",
"10010111000100000101010",
"10010110111100000010111",
"10010110110100000001000",
"10010110101011111111100",
"10010110100011111110101",
"10010110011011111110001",
"10010110010011111110001",
"10010110001011111110101",
"10010110000011111111100",
"10010101111100000001000",
"10010101110100000010111",
"10010101101100000101010",
"10010101100100001000000",
"10010101011100001011011",
"10010101010100001111001",
"10010101001100010011011",
"10010101000100011000000",
"10010100111100011101001",
"10010100110100100010110",
"10010100101100101000111",
"10010100100100101111010",
"10010100011100110110011",
"10010100010100111101110",
"10010100001101000101110",
"10010100000101001110001",
"10010011111101010111000",
"10010011110101100000011",
"10010011101101101010000",
"10010011100101110100010",
"10010011011101111111000",
"10010011010110001010001",
"10010011001110010101101",
"10010011000110100001110",
"10010010111110101110010",
"10010010110110111011001",
"10010010101111001000101",
"10010010100111010110100",
"10010010011111100100110",
"10010010010111110011100",
"10010010010000000010101",
"10010010001000010010011",
"10010010000000100010100",
"10010001111000110011001",
"10010001110001000100000",
"10010001101001010101011",
"10010001100001100111011",
"10010001011001111001110",
"10010001010010001100100",
"10010001001010011111101",
"10010001000010110011011",
"10010000111011000111100",
"10010000110011011100000",
"10010000101011110001000",
"10010000100100000110100",
"10010000011100011100011",
"10010000010100110010101",
"10010000001101001001011",
"10010000000101100000100",
"10001111111101111000001",
"10001111110110010000010",
"10001111101110101000110",
"10001111100111000001101",
"10001111011111011011000",
"10001111010111110100110",
"10001111010000001111000",
"10001111001000101001101",
"10001111000001000100111",
"10001110111001100000010",
"10001110110001111100010",
"10001110101010011000110",
"10001110100010110101100",
"10001110011011010010110",
"10001110010011110000011",
"10001110001100001110100",
"10001110000100101101000",
"10001101111101001100000",
"10001101110101101011011",
"10001101101110001011001",
"10001101100110101011011",
"10001101011111001100001",
"10001101010111101101001",
"10001101010000001110101",
"10001101001000110000100",
"10001101000001010010111",
"10001100111001110101101",
"10001100110010011000110",
"10001100101010111100011",
"10001100100011100000011",
"10001100011100000100110",
"10001100010100101001101",
"10001100001101001111000",
"10001100000101110100101",
"10001011111110011010110",
"10001011110111000001010",
"10001011101111101000010",
"10001011101000001111101",
"10001011100000110111011",
"10001011011001011111100",
"10001011010010001000001",
"10001011001010110001001",
"10001011000011011010100",
"10001010111100000100010",
"10001010110100101110100",
"10001010101101011001001",
"10001010100110000100010",
"10001010011110101111101",
"10001010010111011011100",
"10001010010000000111110",
"10001010001000110100100",
"10001010000001100001100",
"10001001111010001110111",
"10001001110010111100111",
"10001001101011101011010",
"10001001100100011001111",
"10001001011101001001000",
"10001001010101111000011",
"10001001001110101000011",
"10001001000111011000101",
"10001001000000001001010",
"10001000111000111010100",
"10001000110001101100000",
"10001000101010011101110",
"10001000100011010000001",
"10001000011100000010111",
"10001000010100110101111",
"10001000001101101001011",
"10001000000110011101010",
"10000111111111010001101",
"10000111111000000110010",
"10000111110000111011011",
"10000111101001110000110",
"10000111100010100110101",
"10000111011011011100110",
"10000111010100010011011",
"10000111001101001010100",
"10000111000110000001111",
"10000110111110111001110",
"10000110110111110001111",
"10000110110000101010100",
"10000110101001100011100",
"10000110100010011100110",
"10000110011011010110101",
"10000110010100010000110",
"10000110001101001011011",
"10000110000110000110001",
"10000101111111000001100",
"10000101110111111101010",
"10000101110000111001010",
"10000101101001110101101",
"10000101100010110010100",
"10000101011011101111110",
"10000101010100101101011",
"10000101001101101011001",
"10000101000110101001101",
"10000100111111101000011",
"10000100111000100111011",
"10000100110001100111000",
"10000100101010100110111",
"10000100100011100111001",
"10000100011100100111110",
"10000100010101101000110",
"10000100001110101010001",
"10000100000111101011111",
"10000100000000101110000",
"10000011111001110000100",
"10000011110010110011011",
"10000011101011110110101",
"10000011100100111010010",
"10000011011101111110010",
"10000011010111000010101",
"10000011010000000111011",
"10000011001001001100100",
"10000011000010010010000",
"10000010111011010111111",
"10000010110100011110000",
"10000010101101100100101",
"10000010100110101011101",
"10000010011111110010111",
"10000010011000111010110",
"10000010010010000010110",
"10000010001011001011001",
"10000010000100010011111",
"10000001111101011101001",
"10000001110110100110101",
"10000001101111110000101",
"10000001101000111010111",
"10000001100010000101011",
"10000001011011010000100",
"10000001010100011011111",
"10000001001101100111100",
"10000001000110110011101",
"10000001000000000000000",
"10000000111001001100110",
"10000000110010011001111",
"10000000101011100111100",
"10000000100100110101011",
"10000000011110000011100",
"10000000010111010010010",
"10000000010000100001010",
"10000000001001110000100",
"10000000000011000000001",
"01111111111100010000001",
"01111111110101100000100",
"01111111101110110001010",
"01111111101000000010010",
"01111111100001010011110",
"01111111011010100101100",
"01111111010011110111110",
"01111111001101001010010",
"01111111000110011101001",
"01111110111111110000010",
"01111110111001000011111",
"01111110110010010111110",
"01111110101011101011111",
"01111110100101000000100",
"01111110011110010101100",
"01111110010111101010111",
"01111110010001000000100",
"01111110001010010110011",
"01111110000011101100110",
"01111101111101000011100",
"01111101110110011010100",
"01111101101111110010000",
"01111101101001001001101",
"01111101100010100001111",
"01111101011011111010010",
"01111101010101010011000",
"01111101001110101100000",
"01111101001000000101100",
"01111101000001011111010",
"01111100111010111001100",
"01111100110100010100000",
"01111100101101101110110",
"01111100100111001001111",
"01111100100000100101100",
"01111100011010000001010",
"01111100010011011101100",
"01111100001100111010000",
"01111100000110010110111",
"01111011111111110100001",
"01111011111001010001101",
"01111011110010101111100",
"01111011101100001101101",
"01111011100101101100010",
"01111011011111001011001",
"01111011011000101010010",
"01111011010010001001111",
"01111011001011101001110",
"01111011000101001010000",
"01111010111110101010101",
"01111010111000001011100",
"01111010110001101100110",
"01111010101011001110010",
"01111010100100110000001",
"01111010011110010010011",
"01111010010111110100111",
"01111010010001010111111",
"01111010001010111011000",
"01111010000100011110100",
"01111001111110000010100",
"01111001110111100110100",
"01111001110001001011001",
"01111001101010110000000",
"01111001100100010101001",
"01111001011101111010110",
"01111001010111100000101",
"01111001010001000110101",
"01111001001010101101001",
"01111001000100010100000",
"01111000111101111011001",
"01111000110111100010101",
"01111000110001001010011",
"01111000101010110010100",
"01111000100100011011000",
"01111000011110000011110",
"01111000010111101100110",
"01111000010001010110010",
"01111000001010111111111",
"01111000000100101010000",
"01110111111110010100011",
"01110111110111111111000",
"01110111110001101010000",
"01110111101011010101011",
"01110111100101000001000",
"01110111011110101101000",
"01110111011000011001010",
"01110111010010000101111",
"01110111001011110010110",
"01110111000101100000000",
"01110110111111001101100",
"01110110111000111011011",
"01110110110010101001101",
"01110110101100011000000",
"01110110100110000110111",
"01110110011111110110001",
"01110110011001100101100",
"01110110010011010101001",
"01110110001101000101010",
"01110110000110110101101",
"01110110000000100110010",
"01110101111010010111011",
"01110101110100001000101",
"01110101101101111010011",
"01110101100111101100001",
"01110101100001011110100",
"01110101011011010001000",
"01110101010101000011111",
"01110101001110110111001",
"01110101001000101010100",
"01110101000010011110011",
"01110100111100010010100",
"01110100110110000110110",
"01110100101111111011101",
"01110100101001110000101",
"01110100100011100110000",
"01110100011101011011101",
"01110100010111010001100",
"01110100010001000111110",
"01110100001010111110011",
"01110100000100110101001",
"01110011111110101100011",
"01110011111000100011110",
"01110011110010011011101",
"01110011101100010011101",
"01110011100110001100001",
"01110011100000000100101",
"01110011011001111101110",
"01110011010011110111000",
"01110011001101110000101",
"01110011000111101010011",
"01110011000001100100101",
"01110010111011011111001",
"01110010110101011001111",
"01110010101111010101000",
"01110010101001010000010",
"01110010100011001011111",
"01110010011101000111111",
"01110010010111000100010",
"01110010010001000000110",
"01110010001010111101101",
"01110010000100111010111",
"01110001111110111000010",
"01110001111000110110000",
"01110001110010110100000",
"01110001101100110010011",
"01110001100110110001000",
"01110001100000110000000",
"01110001011010101111010",
"01110001010100101110110",
"01110001001110101110100",
"01110001001000101110101",
"01110001000010101111000",
"01110000111100101111110",
"01110000110110110000101",
"01110000110000110010000",
"01110000101010110011100",
"01110000100100110101011",
"01110000011110110111100",
"01110000011000111001111",
"01110000010010111100101",
"01110000001100111111101",
"01110000000111000010111",
"01110000000001000110100",
"01101111111011001010011",
"01101111110101001110100",
"01101111101111010011000",
"01101111101001010111101",
"01101111100011011100110",
"01101111011101100010000",
"01101111010111100111101",
"01101111010001101101101",
"01101111001011110011110",
"01101111000101111010001",
"01101111000000000000111",
"01101110111010000111111",
"01101110110100001111010",
"01101110101110010110110",
"01101110101000011110101",
"01101110100010100110110",
"01101110011100101111001",
"01101110010110110111111",
"01101110010001000000111",
"01101110001011001010001",
"01101110000101010011110",
"01101101111111011101101",
"01101101111001100111101",
"01101101110011110010000",
"01101101101101111100110",
"01101101101000000111110",
"01101101100010010010111",
"01101101011100011110011",
"01101101010110101010001",
"01101101010000110110010",
"01101101001011000010101",
"01101101000101001111010",
"01101100111111011100000",
"01101100111001101001010",
"01101100110011110110110",
"01101100101110000100011",
"01101100101000010010100",
"01101100100010100000110",
"01101100011100101111010",
"01101100010110111110001",
"01101100010001001101001",
"01101100001011011100100",
"01101100000101101100001",
"01101011111111111100001",
"01101011111010001100010",
"01101011110100011100101",
"01101011101110101101011",
"01101011101000111110100",
"01101011100011001111110",
"01101011011101100001010",
"01101011010111110011001",
"01101011010010000101001",
"01101011001100010111100",
"01101011000110101010001",
"01101011000000111101000",
"01101010111011010000010",
"01101010110101100011101",
"01101010101111110111010",
"01101010101010001011010",
"01101010100100011111100",
"01101010011110110100000",
"01101010011001001000110",
"01101010010011011101110",
"01101010001101110011000",
"01101010001000001000101",
"01101010000010011110100",
"01101001110111001010111",
"01101001101011111000011",
"01101001100000100111000",
"01101001010101010110101",
"01101001001010000111010",
"01101000111110111001000",
"01101000110011101011110",
"01101000101000011111100",
"01101000011101010100011",
"01101000010010001010010",
"01101000000111000001001",
"01100111111011111001001",
"01100111110000110010001",
"01100111100101101100001",
"01100111011010100111010",
"01100111001111100011010",
"01100111000100100000011",
"01100110111001011110011",
"01100110101110011101100",
"01100110100011011101101",
"01100110011000011110110",
"01100110001101100001000",
"01100110000010100100001",
"01100101110111101000001",
"01100101101100101101011",
"01100101100001110011100",
"01100101010110111010101",
"01100101001100000010110",
"01100101000001001100000",
"01100100110110010110001",
"01100100101011100001010",
"01100100100000101101010",
"01100100010101111010010",
"01100100001011001000011",
"01100100000000010111100",
"01100011110101100111011",
"01100011101010111000011",
"01100011100000001010011",
"01100011010101011101010",
"01100011001010110001010",
"01100011000000000110000",
"01100010110101011011111",
"01100010101010110010101",
"01100010100000001010010",
"01100010010101100011000",
"01100010001010111100110",
"01100010000000010111010",
"01100001110101110010110",
"01100001101011001111010",
"01100001100000101100101",
"01100001010110001011000",
"01100001001011101010011",
"01100001000001001010100",
"01100000110110101011110",
"01100000101100001101111",
"01100000100001110000111",
"01100000010111010100111",
"01100000001100111001110",
"01100000000010011111100",
"01011111111000000110010",
"01011111101101101101111",
"01011111100011010110100",
"01011111011001000000001",
"01011111001110101010100",
"01011111000100010101110",
"01011110111010000010000",
"01011110101111101111001",
"01011110100101011101010",
"01011110011011001100001",
"01011110010000111100000",
"01011110000110101100101",
"01011101111100011110011",
"01011101110010010000111",
"01011101101000000100011",
"01011101011101111000101",
"01011101010011101101111",
"01011101001001100011111",
"01011100111111011010111",
"01011100110101010010110",
"01011100101011001011100",
"01011100100001000101001",
"01011100010110111111101",
"01011100001100111011000",
"01011100000010110111010",
"01011011111000110100011",
"01011011101110110010011",
"01011011100100110001001",
"01011011011010110000111",
"01011011010000110001100",
"01011011000110110011000",
"01011010111100110101010",
"01011010110010111000100",
"01011010101000111100011",
"01011010011111000001010",
"01011010010101000111000",
"01011010001011001101101",
"01011010000001010101000",
"01011001110111011101010",
"01011001101101100110011",
"01011001100011110000010",
"01011001011001111011001",
"01011001010000000110110",
"01011001000110010011001",
"01011000111100100000100",
"01011000110010101110101",
"01011000101000111101101",
"01011000011111001101011",
"01011000010101011110000",
"01011000001011101111100",
"01011000000010000001110",
"01010111111000010100111",
"01010111101110101000110",
"01010111100100111101100",
"01010111011011010011000",
"01010111010001101001011",
"01010111001000000000101",
"01010110111110011000100",
"01010110110100110001011",
"01010110101011001011000",
"01010110100001100101011",
"01010110011000000000100",
"01010110001110011100100",
"01010110000100111001011",
"01010101111011010110111",
"01010101110001110101011",
"01010101101000010100101",
"01010101011110110100101",
"01010101010101010101011",
"01010101001011110111000",
"01010101000010011001010",
"01010100111000111100100",
"01010100101111100000100",
"01010100100110000101001",
"01010100011100101010101",
"01010100010011010001000",
"01010100001001111000000",
"01010100000000011111111",
"01010011110111001000100",
"01010011101101110001110",
"01010011100100011100000",
"01010011011011000110111",
"01010011010001110010101",
"01010011001000011111001",
"01010010111111001100010",
"01010010110101111010011",
"01010010101100101001000",
"01010010100011011000100",
"01010010011010001000111",
"01010010010000111001111",
"01010010000111101011101",
"01010001111110011110001",
"01010001110101010001100",
"01010001101100000101101",
"01010001100010111010011",
"01010001011001101111111",
"01010001010000100110001",
"01010001000111011101001",
"01010000111110010100111",
"01010000110101001101100",
"01010000101100000110110",
"01010000100011000000110",
"01010000011001111011011",
"01010000010000110110111",
"01010000000111110011001",
"01001111111110110000000",
"01001111110101101101101",
"01001111101100101100000",
"01001111100011101011001",
"01001111011010101011000",
"01001111010001101011101",
"01001111001000101100110",
"01001110111111101110110",
"01001110110110110001100",
"01001110101101110101000",
"01001110100100111001001",
"01001110011011111110000",
"01001110010011000011101",
"01001110001010001001111",
"01001110000001010000111",
"01001101111000011000101",
"01001101101111100001000",
"01001101100110101010001",
"01001101011101110100000",
"01001101010100111110100",
"01001101001100001001110",
"01001101000011010101101",
"01001100111010100010011",
"01001100110001101111101",
"01001100101000111101110",
"01001100100000001100100",
"01001100010111011011111",
"01001100001110101100000",
"01001100000101111100110",
"01001011111101001110010",
"01001011110100100000011",
"01001011101011110011010",
"01001011100011000110111",
"01001011011010011011000",
"01001011010001110000000",
"01001011001001000101100",
"01001011000000011011111",
"01001010110111110010110",
"01001010101111001010011",
"01001010100110100010110",
"01001010011101111011101",
"01001010010101010101011",
"01001010001100101111101",
"01001010000100001010101",
"01001001111011100110010",
"01001001110011000010100",
"01001001101010011111101",
"01001001100001111101010",
"01001001011001011011101",
"01001001010000111010100",
"01001001001000011010001",
"01001000111111111010011",
"01001000110111011011011",
"01001000101110111101000",
"01001000100110011111010",
"01001000011110000010001",
"01001000010101100101110",
"01001000001101001010000",
"01001000000100101110110",
"01000111111100010100011",
"01000111110011111010100",
"01000111101011100001010",
"01000111100011001000110",
"01000111011010110000111",
"01000111010010011001101",
"01000111001010000010111",
"01000111000001101101000",
"01000110111001010111101",
"01000110110001000010111",
"01000110101000101110111",
"01000110100000011011011",
"01000110011000001000101",
"01000110001111110110100",
"01000110000111100100111",
"01000101111111010100000",
"01000101110111000011101",
"01000101101110110100000",
"01000101100110100101000",
"01000101011110010110100",
"01000101010110001000110",
"01000101001101111011101",
"01000101000101101111001",
"01000100111101100011001",
"01000100110101010111111",
"01000100101101001101001",
"01000100100101000011000",
"01000100011100111001101",
"01000100010100110000110",
"01000100001100101000100",
"01000100000100100000111",
"01000011111100011001110",
"01000011110100010011011",
"01000011101100001101101",
"01000011100100001000011",
"01000011011100000011110",
"01000011010011111111110",
"01000011001011111100011",
"01000011000011111001101",
"01000010111011110111100",
"01000010110011110101111",
"01000010101011110100111",
"01000010100011110100100",
"01000010011011110100101",
"01000010010011110101100",
"01000010001011110111000",
"01000010000011111000111",
"01000001111011111011100",
"01000001110011111110101",
"01000001101100000010011",
"01000001100100000110110",
"01000001011100001011101",
"01000001010100010001001",
"01000001001100010111010",
"01000001000100011101111",
"01000000111100100101001",
"01000000110100101101000",
"01000000101100110101100",
"01000000100100111110100",
"01000000011101001000000",
"01000000010101010010001",
"01000000001101011100111",
"01000000000101101000001",
"00111111111101110100001",
"00111111110110000000100",
"00111111101110001101100",
"00111111100110011011001",
"00111111011110101001010",
"00111111010110111000000",
"00111111001111000111010",
"00111111000111010111001",
"00111110111111100111101",
"00111110110111111000101",
"00111110110000001010001",
"00111110101000011100010",
"00111110100000101110110",
"00111110011001000010000",
"00111110010001010101111",
"00111110001001101010001",
"00111110000001111111001",
"00111101111010010100100",
"00111101110010101010100",
"00111101101011000001001",
"00111101100011011000001",
"00111101011011101111111",
"00111101010100001000000",
"00111101001100100000110",
"00111101000100111010001",
"00111100111101010100000",
"00111100110101101110011",
"00111100101110001001011",
"00111100100110100100110",
"00111100011111000000111",
"00111100010111011101011",
"00111100001111111010100",
"00111100001000011000001",
"00111100000000110110011",
"00111011111001010101001",
"00111011110001110100011",
"00111011101010010100001",
"00111011100010110100100",
"00111011011011010101010",
"00111011010011110110101",
"00111011001100011000101",
"00111011000100111011001",
"00111010111101011110001",
"00111010110110000001101",
"00111010101110100101101",
"00111010100111001010010",
"00111010011111101111010",
"00111010011000010100111",
"00111010010000111011001",
"00111010001001100001110",
"00111010000010001000111",
"00111001111010110000101",
"00111001110011011000111",
"00111001101100000001101",
"00111001100100101010111",
"00111001011101010100110",
"00111001010101111111000",
"00111001001110101001111",
"00111001000111010101001",
"00111001000000000001000",
"00111000111000101101011",
"00111000110001011010010",
"00111000101010000111100",
"00111000100010110101100",
"00111000011011100011111",
"00111000010100010010110",
"00111000001101000010010",
"00111000000101110010000",
"00110111111110100010100",
"00110111110111010011011",
"00110111110000000100111",
"00110111101000110110110",
"00110111100001101001010",
"00110111011010011100001",
"00110111010011001111101",
"00110111001100000011100",
"00110111000100110111111",
"00110110111101101100111",
"00110110110110100010010",
"00110110101111011000010",
"00110110101000001110101",
"00110110100001000101100",
"00110110011001111100111",
"00110110010010110100110",
"00110110001011101101001",
"00110110000100100110000",
"00110101111101011111011",
"00110101110110011001010",
"00110101101111010011101",
"00110101101000001110011",
"00110101100001001001101",
"00110101011010000101100",
"00110101010011000001101",
"00110101001011111110011",
"00110101000100111011101",
"00110100111101111001011",
"00110100110110110111100",
"00110100101111110110010",
"00110100101000110101011",
"00110100100001110101000",
"00110100011010110101010",
"00110100010011110101110",
"00110100001100110110111",
"00110100000101111000010",
"00110011111110111010011",
"00110011110111111100111",
"00110011110000111111110",
"00110011101010000011001",
"00110011100011000111001",
"00110011011100001011100",
"00110011010101010000010",
"00110011001110010101100",
"00110011000111011011010",
"00110011000000100001100",
"00110010111001101000010",
"00110010110010101111011",
"00110010101011110111000",
"00110010100100111111001",
"00110010011110000111101",
"00110010010111010000101",
"00110010010000011010001",
"00110010001001100100000",
"00110010000010101110011",
"00110001111011111001010",
"00110001110101000100100",
"00110001101110010000011",
"00110001100111011100100",
"00110001100000101001010",
"00110001011001110110011",
"00110001010011000011111",
"00110001001100010001111",
"00110001000101100000011",
"00110000111110101111010",
"00110000110111111110101",
"00110000110001001110100",
"00110000101010011110110",
"00110000100011101111100",
"00110000011101000000101",
"00110000010110010010011",
"00110000001111100100011",
"00110000001000110110111",
"00110000000010001001110",
"00101111111011011101010",
"00101111110100110001000",
"00101111101110000101010",
"00101111100111011010000",
"00101111100000101111010",
"00101111011010000100110",
"00101111010011011010111",
"00101111001100110001010",
"00101111000110001000001",
"00101110111111011111100",
"00101110111000110111010",
"00101110110010001111100",
"00101110101011101000001",
"00101110100101000001010",
"00101110011110011010110",
"00101110010111110100110",
"00101110010001001111001",
"00101110001010101001111",
"00101110000100000101001",
"00101101111101100000110",
"00101101110110111100111",
"00101101110000011001011",
"00101101101001110110011",
"00101101100011010011110",
"00101101011100110001100",
"00101101010110001111110",
"00101101001111101110011",
"00101101001001001101100",
"00101101000010101101000",
"00101100111100001100111",
"00101100110101101101010",
"00101100101111001110000",
"00101100101000101111001",
"00101100100010010000110",
"00101100011011110010110",
"00101100010101010101001",
"00101100001110111000001",
"00101100001000011011011",
"00101100000001111111000",
"00101011111011100011001",
"00101011110101000111101",
"00101011101110101100100",
"00101011101000010001110",
"00101011100001110111101",
"00101011011011011101110",
"00101011010101000100010",
"00101011001110101011010",
"00101011001000010010101",
"00101011000001111010100",
"00101010111011100010101",
"00101010110101001011010",
"00101010101110110100010",
"00101010101000011101110",
"00101010100010000111100",
"00101010011011110001110",
"00101010010101011100011",
"00101010001111000111011",
"00101010001000110010111",
"00101010000010011110101",
"00101001111100001011000",
"00101001110101110111100",
"00101001101111100100101",
"00101001101001010010000",
"00101001100010111111111",
"00101001011100101110001",
"00101001010110011100110",
"00101001010000001011110",
"00101001001001111011010",
"00101001000011101011000",
"00101000111101011011010",
"00101000110111001011111",
"00101000110000111100111",
"00101000101010101110010",
"00101000100100100000000",
"00101000011110010010001",
"00101000011000000100110",
"00101000010001110111110",
"00101000001011101011001",
"00101000000101011110110",
"00100111111111010011000",
"00100111111001000111100",
"00100111110010111100011",
"00100111101100110001101",
"00100111100110100111010",
"00100111100000011101011",
"00100111011010010011111",
"00100111010100001010101",
"00100111001110000001111",
"00100111000111111001011",
"00100111000001110001011",
"00100110111011101001110",
"00100110110101100010100",
"00100110101111011011100",
"00100110101001010101000",
"00100110100011001111000",
"00100110011101001001010",
"00100110010111000011110",
"00100110010000111110110",
"00100110001010111010010",
"00100110000100110110000",
"00100101111110110010000",
"00100101111000101110100",
"00100101110010101011100",
"00100101101100101000110",
"00100101100110100110010",
"00100101100000100100011",
"00100101011010100010101",
"00100101010100100001011",
"00100101001110100000100",
"00100101001000100000000",
"00100101000010011111111",
"00100100111100100000001",
"00100100110110100000101",
"00100100110000100001100",
"00100100101010100010111",
"00100100100100100100101",
"00100100011110100110101",
"00100100011000101001001",
"00100100010010101011110",
"00100100001100101111000",
"00100100000110110010100",
"00100100000000110110011",
"00100011111010111010101",
"00100011110100111111010",
"00100011101111000100001",
"00100011101001001001011",
"00100011100011001111001",
"00100011011101010101001",
"00100011010111011011100",
"00100011010001100010010",
"00100011001011101001011",
"00100011000101110000111",
"00100010111111111000101",
"00100010111010000000111",
"00100010110100001001011",
"00100010101110010010010",
"00100010101000011011100",
"00100010100010100101001",
"00100010011100101111000",
"00100010010110111001010",
"00100010010001000100000",
"00100010001011001111000",
"00100010000101011010011",
"00100001111111100110000",
"00100001111001110010001",
"00100001110011111110100",
"00100001101110001011010",
"00100001101000011000011",
"00100001100010100101110",
"00100001011100110011101",
"00100001010111000001110",
"00100001010001010000001",
"00100001001011011111000",
"00100001000101101110010",
"00100000111111111101110",
"00100000111010001101101",
"00100000110100011101111",
"00100000101110101110011",
"00100000101000111111010",
"00100000100011010000100",
"00100000011101100010001",
"00100000010111110100000",
"00100000010010000110010",
"00100000001100011000111",
"00100000000110101011110",
"00100000000000111111000",
"00011111111011010010101",
"00011111110101100110101",
"00011111101111111010111",
"00011111101010001111100",
"00011111100100100100011",
"00011111011110111001110",
"00011111011001001111011",
"00011111010011100101010",
"00011111001101111011101",
"00011111001000010010010",
"00011111000010101001010",
"00011110111101000000100",
"00011110110111011000001",
"00011110110001110000001",
"00011110101100001000011",
"00011110100110100001000",
"00011110100000111001111",
"00011110011011010011010",
"00011110010101101100111",
"00011110010000000110110",
"00011110001010100001000",
"00011110000100111011101",
"00011101111111010110100",
"00011101111001110001110",
"00011101110100001101011",
"00011101101110101001010",
"00011101101001000101100",
"00011101100011100010000",
"00011101011101111110111",
"00011101011000011100000",
"00011101010010111001101",
"00011101001101010111011",
"00011101000111110101100",
"00011101000010010100000",
"00011100111100110010111",
"00011100110111010010000",
"00011100110001110001011",
"00011100101100010001001",
"00011100100110110001010",
"00011100100001010001101",
"00011100011011110010011",
"00011100010110010011011",
"00011100010000110100110",
"00011100001011010110011",
"00011100000101111000011",
"00011100000000011010101",
"00011011111010111101010",
"00011011110101100000010",
"00011011110000000011011",
"00011011101010100111000",
"00011011100101001010111",
"00011011011111101111000",
"00011011011010010011100",
"00011011010100111000011",
"00011011001111011101011",
"00011011001010000010111",
"00011011000100101000101",
"00011010111111001110101",
"00011010111001110101000",
"00011010110100011011101",
"00011010101111000010101",
"00011010101001101001111",
"00011010100100010001100",
"00011010011110111001011",
"00011010011001100001101",
"00011010010100001010001",
"00011010001110110010111",
"00011010001001011100000",
"00011010000100000101100",
"00011001111110101111010",
"00011001111001011001010",
"00011001110100000011100",
"00011001101110101110010",
"00011001101001011001001",
"00011001100100000100011",
"00011001011110110000000",
"00011001011001011011110",
"00011001010100000111111",
"00011001001110110100011",
"00011001001001100001001",
"00011001000100001110010",
"00011000111110111011101",
"00011000111001101001010",
"00011000110100010111001",
"00011000101111000101011",
"00011000101001110011111",
"00011000100100100010110",
"00011000011111010001111",
"00011000011010000001011",
"00011000010100110001000",
"00011000001111100001001",
"00011000001010010001011",
"00011000000101000010000",
"00010111111111110010111",
"00010111111010100100000",
"00010111110101010101100",
"00010111110000000111011",
"00010111101010111001011",
"00010111100101101011110",
"00010111100000011110100",
"00010111011011010001011",
"00010111010110000100101",
"00010111010000111000001",
"00010111001011101100000",
"00010111000110100000001",
"00010111000001010100100",
"00010110111100001001010",
"00010110110110111110001",
"00010110110001110011011",
"00010110101100101001000",
"00010110100111011110111",
"00010110100010010101000",
"00010110011101001011011",
"00010110011000000010000",
"00010110010010111001000",
"00010110001101110000011",
"00010110001000100111111",
"00010110000011011111101",
"00010101111110010111110",
"00010101111001010000001",
"00010101110100001000111",
"00010101101111000001110",
"00010101101001111011001",
"00010101100100110100101",
"00010101011111101110011",
"00010101011010101000100",
"00010101010101100010111",
"00010101010000011101100",
"00010101001011011000011",
"00010101000110010011101",
"00010101000001001111001",
"00010100111100001010111",
"00010100110111000110111",
"00010100110010000011001",
"00010100101100111111111",
"00010100100111111100101",
"00010100100010111001111",
"00010100011101110111010",
"00010100011000110101000",
"00010100010011110010111",
"00010100001110110001001",
"00010100001001101111110",
"00010100000100101110100",
"00010011111111101101100",
"00010011111010101100111",
"00010011110101101100100",
"00010011110000101100011",
"00010011101011101100101",
"00010011100110101101000",
"00010011100001101101101",
"00010011011100101110110",
"00010011010111101111111",
"00010011010010110001100",
"00010011001101110011010",
"00010011001000110101010",
"00010011000011110111101",
"00010010111110111010010",
"00010010111001111101000",
"00010010110101000000001",
"00010010110000000011100",
"00010010101011000111010",
"00010010100110001011001",
"00010010100001001111011",
"00010010011100010011110",
"00010010010111011000100",
"00010010010010011101100",
"00010010001101100010110",
"00010010001000101000010",
"00010010000011101110000",
"00010001111110110100001",
"00010001111001111010100",
"00010001110101000001000",
"00010001110000000111110",
"00010001101011001111000",
"00010001100110010110010",
"00010001100001011101111",
"00010001011100100101110",
"00010001010111101101111",
"00010001010010110110011",
"00010001001101111111000",
"00010001001001000111111",
"00010001000100010001001",
"00010000111111011010100",
"00010000111010100100010",
"00010000110101101110001",
"00010000110000111000011",
"00010000101100000010111",
"00010000100111001101101",
"00010000100010011000100",
"00010000011101100011110",
"00010000011000101111011",
"00010000010011111011001",
"00010000001111000111001",
"00010000001010010011011",
"00010000000101011111111",
"00010000000000101100101",
"00001111111011111001101",
"00001111110111000111000",
"00001111110010010100100",
"00001111101101100010010",
"00001111101000110000011",
"00001111100011111110101",
"00001111011111001101001",
"00001111011010011100000",
"00001111010101101011000",
"00001111010000111010010",
"00001111001100001001111",
"00001111000111011001101",
"00001111000010101001110",
"00001110111101111010000",
"00001110111001001010100",
"00001110110100011011011",
"00001110101111101100011",
"00001110101010111101101",
"00001110100110001111010",
"00001110100001100001000",
"00001110011100110011000",
"00001110011000000101011",
"00001110010011010111111",
"00001110001110101010101",
"00001110001001111101101",
"00001110000101010000111",
"00001110000000100100011",
"00001101111011111000001",
"00001101110111001100001",
"00001101110010100000011",
"00001101101101110100111",
"00001101101001001001101",
"00001101100100011110100",
"00001101011111110011110",
"00001101011011001001010",
"00001101010110011110111",
"00001101010001110100111",
"00001101001101001011000",
"00001101001000100001100",
"00001101000011111000001",
"00001100111111001111001",
"00001100111010100110001",
"00001100110101111101101",
"00001100110001010101010",
"00001100101100101101001",
"00001100101000000101001",
"00001100100011011101100",
"00001100011110110110001",
"00001100011010001110111",
"00001100010101101000000",
"00001100010001000001010",
"00001100001100011010111",
"00001100000111110100100",
"00001100000011001110101",
"00001011111110101000111",
"00001011111010000011011",
"00001011110101011110000",
"00001011110000111001000",
"00001011101100010100001",
"00001011100111101111100",
"00001011100011001011001",
"00001011011110100111000",
"00001011011010000011001",
"00001011010101011111100",
"00001011010000111100001",
"00001011001100011001000",
"00001011000111110110000",
"00001011000011010011010",
"00001010111110110000110",
"00001010111010001110100",
"00001010110101101100100",
"00001010110001001010101",
"00001010101100101001001",
"00001010101000000111110",
"00001010100011100110101",
"00001010011111000101110",
"00001010011010100101001",
"00001010010110000100110",
"00001010010001100100100",
"00001010001101000100100",
"00001010001000100100110",
"00001010000100000101011",
"00001001111111100110000",
"00001001111011000111000",
"00001001110110101000001",
"00001001110010001001100",
"00001001101101101011001",
"00001001101001001101000",
"00001001100100101111001",
"00001001100000010001011",
"00001001011011110011111",
"00001001010111010110110",
"00001001010010111001101",
"00001001001110011100111",
"00001001001010000000010",
"00001001000101100011111",
"00001001000001000111110",
"00001000111100101011111",
"00001000111000010000010",
"00001000110011110100110",
"00001000101111011001100",
"00001000101010111110100",
"00001000100110100011110",
"00001000100010001001001",
"00001000011101101110111",
"00001000011001010100101",
"00001000010100111010110",
"00001000010000100001000",
"00001000001100000111101",
"00001000000111101110011",
"00001000000011010101010",
"00000111111110111100100",
"00000111111010100011111",
"00000111110110001011100",
"00000111110001110011011",
"00000111101101011011011",
"00000111101001000011110",
"00000111100100101100001",
"00000111100000010100111",
"00000111011011111101111",
"00000111010111100110111",
"00000111010011010000011",
"00000111001110111001111",
"00000111001010100011101",
"00000111000110001101101",
"00000111000001110111111",
"00000110111101100010010",
"00000110111001001101000",
"00000110110100110111111",
"00000110110000100010111",
"00000110101100001110001",
"00000110100111111001110",
"00000110100011100101100",
"00000110011111010001011",
"00000110011010111101100",
"00000110010110101001111",
"00000110010010010110100",
"00000110001110000011010",
"00000110001001110000010",
"00000110000101011101011",
"00000110000001001010111",
"00000101111100111000011",
"00000101111000100110010",
"00000101110100010100011",
"00000101110000000010100",
"00000101101011110001000",
"00000101100111011111101",
"00000101100011001110101",
"00000101011110111101110",
"00000101011010101101000",
"00000101010110011100100",
"00000101010010001100001",
"00000101001101111100001",
"00000101001001101100010",
"00000101000101011100100",
"00000101000001001101001",
"00000100111100111101111",
"00000100111000101110111",
"00000100110100100000000",
"00000100110000010001011",
"00000100101100000010111",
"00000100100111110100110",
"00000100100011100110101",
"00000100011111011000111",
"00000100011011001011010",
"00000100010110111101111",
"00000100010010110000101",
"00000100001110100011101",
"00000100001010010110111",
"00000100000110001010010",
"00000100000001111101111",
"00000011111101110001110",
"00000011111001100101110",
"00000011110101011010000",
"00000011110001001110011",
"00000011101101000011000",
"00000011101000110111111",
"00000011100100101100111",
"00000011100000100010001",
"00000011011100010111100",
"00000011011000001101001",
"00000011010100000011000",
"00000011001111111001000",
"00000011001011101111010",
"00000011000111100101101",
"00000011000011011100011",
"00000010111111010011001",
"00000010111011001010001",
"00000010110111000001011",
"00000010110010111000111",
"00000010101110110000100",
"00000010101010101000010",
"00000010100110100000010",
"00000010100010011000100",
"00000010011110010000111",
"00000010011010001001100",
"00000010010110000010011",
"00000010010001111011011",
"00000010001101110100100",
"00000010001001101101111",
"00000010000101100111100",
"00000010000001100001010",
"00000001111101011011010",
"00000001111001010101100",
"00000001110101001111111",
"00000001110001001010011",
"00000001101101000101001",
"00000001101001000000000",
"00000001100100111011010",
"00000001100000110110100",
"00000001011100110010001",
"00000001011000101101111",
"00000001010100101001110",
"00000001010000100101110",
"00000001001100100010001",
"00000001001000011110101",
"00000001000100011011010",
"00000001000000011000010",
"00000000111100010101010",
"00000000111000010010100",
"00000000110100010000000",
"00000000110000001101100",
"00000000101100001011011",
"00000000101000001001011",
"00000000100100000111101",
"00000000100000000110000",
"00000000011100000100101",
"00000000011000000011011",
"00000000010100000010011",
"00000000010000000001100",
"00000000001100000000111",
"00000000001000000000011",
"00000000000100000000001");

begin

  data<=rom1(conv_integer(addr));
  data2<=rom2(conv_integer(addr));

  end VHDL;
