/home/mizuta1018/HW/FPU/VHDL/fsin/fmul_3.vhd