library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

entity invromfetch is
  port(addr: in std_logic_vector(10 downto 0);
       data,data2:  out std_logic_vector(22 downto 0) -- 23bit
       );
  end invromfetch;

architecture VHDL of invromfetch is

  type rom_t is array(0 to 2047) of std_logic_vector(22 downto 0);
  constant rom1 : rom_t :=("11111111111111111111111",
"11111111110000000000100",
"11111111100000000010000",
"11111111010000000100100",
"11111111000000001000000",
"11111110110000001100100",
"11111110100000010010000",
"11111110010000011000100",
"11111110000000100000000",
"11111101110000101000011",
"11111101100000110001111",
"11111101010000111100010",
"11111101000001000111101",
"11111100110001010100000",
"11111100100001100001011",
"11111100010001101111110",
"11111100000001111111001",
"11111011110010001111011",
"11111011100010100000101",
"11111011010010110010111",
"11111011000011000110001",
"11111010110011011010011",
"11111010100011101111100",
"11111010010100000101101",
"11111010000100011100110",
"11111001110100110100110",
"11111001100101001101111",
"11111001010101100111111",
"11111001000110000010110",
"11111000110110011110110",
"11111000100110111011101",
"11111000010111011001011",
"11111000000111111000001",
"11110111111000010111111",
"11110111101000111000101",
"11110111011001011010010",
"11110111001001111100111",
"11110110111010100000011",
"11110110101011000100111",
"11110110011011101010011",
"11110110001100010000110",
"11110101111100111000001",
"11110101101101100000011",
"11110101011110001001100",
"11110101001110110011110",
"11110100111111011110110",
"11110100110000001010111",
"11110100100000110111110",
"11110100010001100101101",
"11110100000010010100100",
"11110011110011000100010",
"11110011100011110101000",
"11110011010100100110101",
"11110011000101011001001",
"11110010110110001100101",
"11110010100111000001000",
"11110010010111110110011",
"11110010001000101100101",
"11110001111001100011110",
"11110001101010011011111",
"11110001011011010100111",
"11110001001100001110110",
"11110000111101001001101",
"11110000101110000101011",
"11110000011111000010000",
"11110000001111111111101",
"11110000000000111110000",
"11101111110001111101100",
"11101111100010111101110",
"11101111010011111111000",
"11101111000101000001001",
"11101110110110000100001",
"11101110100111001000000",
"11101110011000001100111",
"11101110001001010010101",
"11101101111010011001010",
"11101101101011100000110",
"11101101011100101001001",
"11101101001101110010100",
"11101100111110111100101",
"11101100110000000111110",
"11101100100001010011110",
"11101100010010100000101",
"11101100000011101110011",
"11101011110100111101000",
"11101011100110001100101",
"11101011010111011101000",
"11101011001000101110011",
"11101010111010000000100",
"11101010101011010011101",
"11101010011100100111101",
"11101010001101111100011",
"11101001111111010010001",
"11101001110000101000110",
"11101001100010000000001",
"11101001010011011000100",
"11101001000100110001110",
"11101000110110001011111",
"11101000100111100110110",
"11101000011001000010101",
"11101000001010011111010",
"11100111111011111100111",
"11100111101101011011010",
"11100111011110111010100",
"11100111010000011010110",
"11100111000001111011110",
"11100110110011011101101",
"11100110100101000000011",
"11100110010110100011111",
"11100110001000001000011",
"11100101111001101101101",
"11100101101011010011111",
"11100101011100111010111",
"11100101001110100010110",
"11100101000000001011011",
"11100100110001110101000",
"11100100100011011111011",
"11100100010101001010101",
"11100100000110110110110",
"11100011111000100011110",
"11100011101010010001100",
"11100011011100000000001",
"11100011001101101111101",
"11100010111111100000000",
"11100010110001010001001",
"11100010100011000011001",
"11100010010100110110000",
"11100010000110101001101",
"11100001111000011110001",
"11100001101010010011100",
"11100001011100001001110",
"11100001001110000000110",
"11100000111111111000100",
"11100000110001110001010",
"11100000100011101010110",
"11100000010101100101000",
"11100000000111100000001",
"11011111111001011100001",
"11011111101011011001000",
"11011111011101010110100",
"11011111001111010101000",
"11011111000001010100010",
"11011110110011010100011",
"11011110100101010101010",
"11011110010111010111000",
"11011110001001011001100",
"11011101111011011100111",
"11011101101101100001000",
"11011101011111100110000",
"11011101010001101011110",
"11011101000011110010010",
"11011100110101111001110",
"11011100101000000001111",
"11011100011010001010111",
"11011100001100010100110",
"11011011111110011111011",
"11011011110000101010110",
"11011011100010110111000",
"11011011010101000100000",
"11011011000111010001111",
"11011010111001100000100",
"11011010101011110000000",
"11011010011110000000001",
"11011010010000010001010",
"11011010000010100011000",
"11011001110100110101101",
"11011001100111001001000",
"11011001011001011101010",
"11011001001011110010010",
"11011000111110001000000",
"11011000110000011110100",
"11011000100010110101111",
"11011000010101001110000",
"11011000000111100110111",
"11010111111010000000101",
"11010111101100011011001",
"11010111011110110110011",
"11010111010001010010011",
"11010111000011101111010",
"11010110110110001100111",
"11010110101000101011010",
"11010110011011001010011",
"11010110001101101010011",
"11010110000000001011001",
"11010101110010101100100",
"11010101100101001110111",
"11010101010111110001111",
"11010101001010010101101",
"11010100111100111010010",
"11010100101111011111100",
"11010100100010000101101",
"11010100010100101100100",
"11010100000111010100001",
"11010011111001111100101",
"11010011101100100101110",
"11010011011111001111101",
"11010011010001111010011",
"11010011000100100101110",
"11010010110111010010000",
"11010010101001111111000",
"11010010011100101100110",
"11010010001111011011001",
"11010010000010001010011",
"11010001110100111010011",
"11010001100111101011001",
"11010001011010011100101",
"11010001001101001110111",
"11010001000000000001111",
"11010000110010110101101",
"11010000100101101010001",
"11010000011000011111011",
"11010000001011010101011",
"11001111111110001100000",
"11001111110001000011100",
"11001111100011111011110",
"11001111010110110100110",
"11001111001001101110011",
"11001110111100101000111",
"11001110101111100100000",
"11001110100010100000000",
"11001110010101011100101",
"11001110001000011010000",
"11001101111011011000001",
"11001101101110010111000",
"11001101100001010110101",
"11001101010100010110111",
"11001101000111011000000",
"11001100111010011001110",
"11001100101101011100010",
"11001100100000011111100",
"11001100010011100011100",
"11001100000110101000010",
"11001011111001101101101",
"11001011101100110011110",
"11001011011111111010101",
"11001011010011000010010",
"11001011000110001010101",
"11001010111001010011101",
"11001010101100011101011",
"11001010011111100111111",
"11001010010010110011001",
"11001010000101111111000",
"11001001111001001011101",
"11001001101100011001000",
"11001001011111100111000",
"11001001010010110101110",
"11001001000110000101010",
"11001000111001010101100",
"11001000101100100110011",
"11001000011111111000000",
"11001000010011001010011",
"11001000000110011101011",
"11000111111001110001001",
"11000111101101000101101",
"11000111100000011010110",
"11000111010011110000101",
"11000111000111000111001",
"11000110111010011110011",
"11000110101101110110011",
"11000110100001001111000",
"11000110010100101000011",
"11000110001000000010100",
"11000101111011011101010",
"11000101101110111000110",
"11000101100010010100111",
"11000101010101110001110",
"11000101001001001111010",
"11000100111100101101100",
"11000100110000001100011",
"11000100100011101100000",
"11000100010111001100011",
"11000100001010101101011",
"11000011111110001111000",
"11000011110001110001011",
"11000011100101010100100",
"11000011011000111000010",
"11000011001100011100110",
"11000011000000000001110",
"11000010110011100111101",
"11000010100111001110001",
"11000010011010110101010",
"11000010001110011101001",
"11000010000010000101101",
"11000001110101101110111",
"11000001101001011000110",
"11000001011101000011010",
"11000001010000101110100",
"11000001000100011010100",
"11000000111000000111000",
"11000000101011110100011",
"11000000011111100010010",
"11000000010011010000111",
"11000000000111000000001",
"10111111111010110000001",
"10111111101110100000110",
"10111111100010010010000",
"10111111010110000100000",
"10111111001001110110101",
"10111110111101101001111",
"10111110110001011101111",
"10111110100101010010100",
"10111110011001000111110",
"10111110001100111101110",
"10111110000000110100011",
"10111101110100101011101",
"10111101101000100011100",
"10111101011100011100001",
"10111101010000010101011",
"10111101000100001111010",
"10111100111000001001111",
"10111100101100000101000",
"10111100100000000000111",
"10111100010011111101100",
"10111100000111111010101",
"10111011111011111000100",
"10111011101111110111000",
"10111011100011110110001",
"10111011010111110101111",
"10111011001011110110010",
"10111010111111110111011",
"10111010110011111001001",
"10111010100111111011100",
"10111010011011111110100",
"10111010010000000010010",
"10111010000100000110100",
"10111001111000001011100",
"10111001101100010001001",
"10111001100000010111011",
"10111001010100011110010",
"10111001001000100101110",
"10111000111100101101111",
"10111000110000110110110",
"10111000100101000000001",
"10111000011001001010010",
"10111000001101010101000",
"10111000000001100000010",
"10110111110101101100010",
"10110111101001111000111",
"10110111011110000110001",
"10110111010010010100000",
"10110111000110100010101",
"10110110111010110001110",
"10110110101111000001100",
"10110110100011010001111",
"10110110010111100010111",
"10110110001011110100101",
"10110110000000000110111",
"10110101110100011001110",
"10110101101000101101011",
"10110101011101000001100",
"10110101010001010110010",
"10110101000101101011110",
"10110100111010000001110",
"10110100101110011000011",
"10110100100010101111101",
"10110100010111000111101",
"10110100001011100000001",
"10110011111111111001010",
"10110011110100010011000",
"10110011101000101101011",
"10110011011101001000011",
"10110011010001100011111",
"10110011000110000000001",
"10110010111010011101000",
"10110010101110111010011",
"10110010100011011000100",
"10110010010111110111001",
"10110010001100010110011",
"10110010000000110110010",
"10110001110101010110110",
"10110001101001110111111",
"10110001011110011001101",
"10110001010010111011111",
"10110001000111011110111",
"10110000111100000010011",
"10110000110000100110100",
"10110000100101001011010",
"10110000011001110000101",
"10110000001110010110100",
"10110000000010111101001",
"10101111110111100100010",
"10101111101100001100000",
"10101111100000110100010",
"10101111010101011101010",
"10101111001010000110110",
"10101110111110110000111",
"10101110110011011011101",
"10101110101000000111000",
"10101110011100110010111",
"10101110010001011111011",
"10101110000110001100100",
"10101101111010111010010",
"10101101101111101000100",
"10101101100100010111011",
"10101101011001000110111",
"10101101001101110111000",
"10101101000010100111101",
"10101100110111011000111",
"10101100101100001010110",
"10101100100000111101001",
"10101100010101110000001",
"10101100001010100011110",
"10101011111111010111111",
"10101011110100001100101",
"10101011101001000010000",
"10101011011101111000000",
"10101011010010101110100",
"10101011000111100101100",
"10101010111100011101010",
"10101010110001010101100",
"10101010100110001110010",
"10101010011011000111110",
"10101010010000000001110",
"10101010000100111100010",
"10101001111001110111011",
"10101001101110110011001",
"10101001100011101111011",
"10101001011000101100010",
"10101001001101101001110",
"10101001000010100111110",
"10101000110111100110011",
"10101000101100100101100",
"10101000100001100101010",
"10101000010110100101100",
"10101000001011100110011",
"10101000000000100111110",
"10100111110101101001110",
"10100111101010101100011",
"10100111011111101111100",
"10100111010100110011010",
"10100111001001110111100",
"10100110111110111100010",
"10100110110100000001110",
"10100110101001000111101",
"10100110011110001110001",
"10100110010011010101010",
"10100110001000011100111",
"10100101111101100101001",
"10100101110010101101111",
"10100101100111110111010",
"10100101011101000001001",
"10100101010010001011100",
"10100101000111010110100",
"10100100111100100010000",
"10100100110001101110001",
"10100100100110111010111",
"10100100011100001000000",
"10100100010001010101111",
"10100100000110100100001",
"10100011111011110011000",
"10100011110001000010100",
"10100011100110010010011",
"10100011011011100011000",
"10100011010000110100000",
"10100011000110000101101",
"10100010111011010111111",
"10100010110000101010101",
"10100010100101111101111",
"10100010011011010001101",
"10100010010000100110000",
"10100010000101111010111",
"10100001111011010000011",
"10100001110000100110011",
"10100001100101111100111",
"10100001011011010100000",
"10100001010000101011101",
"10100001000110000011110",
"10100000111011011100100",
"10100000110000110101110",
"10100000100110001111100",
"10100000011011101001111",
"10100000010001000100110",
"10100000000110100000001",
"10011111111011111100001",
"10011111110001011000100",
"10011111100110110101101",
"10011111011100010011001",
"10011111010001110001001",
"10011111000111001111110",
"10011110111100101111000",
"10011110110010001110101",
"10011110100111101110111",
"10011110011101001111101",
"10011110010010110000111",
"10011110001000010010101",
"10011101111101110101000",
"10011101110011010111111",
"10011101101000111011010",
"10011101011110011111001",
"10011101010100000011101",
"10011101001001101000100",
"10011100111111001110000",
"10011100110100110100000",
"10011100101010011010101",
"10011100100000000001101",
"10011100010101101001010",
"10011100001011010001011",
"10011100000000111010000",
"10011011110110100011001",
"10011011101100001100110",
"10011011100001110111000",
"10011011010111100001110",
"10011011001101001101000",
"10011011000010111000101",
"10011010111000100101000",
"10011010101110010001110",
"10011010100011111111000",
"10011010011001101100111",
"10011010001111011011001",
"10011010000101001010000",
"10011001111010111001011",
"10011001110000101001010",
"10011001100110011001101",
"10011001011100001010100",
"10011001010001111100000",
"10011001000111101101111",
"10011000111101100000010",
"10011000110011010011010",
"10011000101001000110101",
"10011000011110111010101",
"10011000010100101111001",
"10011000001010100100000",
"10011000000000011001100",
"10010111110110001111100",
"10010111101100000110000",
"10010111100001111101000",
"10010111010111110100100",
"10010111001101101100100",
"10010111000011100101000",
"10010110111001011110000",
"10010110101111010111100",
"10010110100101010001100",
"10010110011011001100000",
"10010110010001000111000",
"10010110000111000010101",
"10010101111100111110101",
"10010101110010111011001",
"10010101101000111000001",
"10010101011110110101101",
"10010101010100110011101",
"10010101001010110010001",
"10010101000000110001001",
"10010100110110110000101",
"10010100101100110000100",
"10010100100010110001000",
"10010100011000110010000",
"10010100001110110011100",
"10010100000100110101011",
"10010011111010110111111",
"10010011110000111010110",
"10010011100110111110010",
"10010011011101000010001",
"10010011010011000110100",
"10010011001001001011011",
"10010010111111010000110",
"10010010110101010110101",
"10010010101011011101000",
"10010010100001100011111",
"10010010010111101011010",
"10010010001101110011000",
"10010010000011111011011",
"10010001111010000100001",
"10010001110000001101011",
"10010001100110010111001",
"10010001011100100001011",
"10010001010010101100001",
"10010001001000110111010",
"10010000111111000011000",
"10010000110101001111001",
"10010000101011011011110",
"10010000100001101000111",
"10010000010111110110100",
"10010000001110000100100",
"10010000000100010011001",
"10001111111010100010001",
"10001111110000110001101",
"10001111100111000001101",
"10001111011101010010000",
"10001111010011100011000",
"10001111001001110100011",
"10001111000000000110010",
"10001110110110011000101",
"10001110101100101011100",
"10001110100010111110110",
"10001110011001010010100",
"10001110001111100110110",
"10001110000101111011100",
"10001101111100010000101",
"10001101110010100110010",
"10001101101000111100011",
"10001101011111010011000",
"10001101010101101010001",
"10001101001100000001101",
"10001101000010011001101",
"10001100111000110010000",
"10001100101111001011000",
"10001100100101100100011",
"10001100011011111110010",
"10001100010010011000100",
"10001100001000110011010",
"10001011111111001110100",
"10001011110101101010010",
"10001011101100000110011",
"10001011100010100011000",
"10001011011001000000001",
"10001011001111011101101",
"10001011000101111011110",
"10001010111100011010001",
"10001010110010111001001",
"10001010101001011000100",
"10001010011111111000011",
"10001010010110011000101",
"10001010001100111001011",
"10001010000011011010101",
"10001001111001111100010",
"10001001110000011110011",
"10001001100111000001000",
"10001001011101100100000",
"10001001010100000111100",
"10001001001010101011100",
"10001001000001001111111",
"10001000110111110100110",
"10001000101110011010000",
"10001000100100111111110",
"10001000011011100110000",
"10001000010010001100101",
"10001000001000110011110",
"10000111111111011011010",
"10000111110110000011010",
"10000111101100101011110",
"10000111100011010100101",
"10000111011001111110000",
"10000111010000100111110",
"10000111000111010010000",
"10000110111101111100110",
"10000110110100100111111",
"10000110101011010011011",
"10000110100001111111011",
"10000110011000101011111",
"10000110001111011000110",
"10000110000110000110001",
"10000101111100110011111",
"10000101110011100010001",
"10000101101010010000111",
"10000101100001000000000",
"10000101010111101111100",
"10000101001110011111100",
"10000101000101001111111",
"10000100111100000000110",
"10000100110010110010001",
"10000100101001100011111",
"10000100100000010110000",
"10000100010111001000101",
"10000100001101111011110",
"10000100000100101111010",
"10000011111011100011001",
"10000011110010010111100",
"10000011101001001100010",
"10000011100000000001100",
"10000011010110110111010",
"10000011001101101101011",
"10000011000100100011111",
"10000010111011011010111",
"10000010110010010010010",
"10000010101001001010000",
"10000010100000000010010",
"10000010010110111011000",
"10000010001101110100001",
"10000010000100101101101",
"10000001111011100111101",
"10000001110010100010000",
"10000001101001011100111",
"10000001100000011000001",
"10000001010111010011111",
"10000001001110001111111",
"10000001000101001100100",
"10000000111100001001011",
"10000000110011000110111",
"10000000101010000100101",
"10000000100001000010111",
"10000000011000000001100",
"10000000001111000000101",
"10000000000110000000001",
"01111111111101000000000",
"01111111110100000000011",
"01111111101011000001001",
"01111111100010000010011",
"01111111011001000100000",
"01111111010000000110000",
"01111111000111001000100",
"01111110111110001011011",
"01111110110101001110101",
"01111110101100010010011",
"01111110100011010110100",
"01111110011010011011000",
"01111110010001100000000",
"01111110001000100101011",
"01111101111111101011001",
"01111101110110110001011",
"01111101101101111000000",
"01111101100100111111000",
"01111101011100000110100",
"01111101010011001110011",
"01111101001010010110101",
"01111101000001011111010",
"01111100111000101000011",
"01111100101111110001111",
"01111100100110111011111",
"01111100011110000110001",
"01111100010101010000111",
"01111100001100011100000",
"01111100000011100111101",
"01111011111010110011101",
"01111011110010000000000",
"01111011101001001100110",
"01111011100000011010000",
"01111011010111100111101",
"01111011001110110101101",
"01111011000110000100000",
"01111010111101010010111",
"01111010110100100010001",
"01111010101011110001110",
"01111010100011000001110",
"01111010011010010010001",
"01111010010001100011000",
"01111010001000110100010",
"01111010000000000101111",
"01111001110111011000000",
"01111001101110101010100",
"01111001100101111101010",
"01111001011101010000101",
"01111001010100100100010",
"01111001001011111000010",
"01111001000011001100110",
"01111000111010100001101",
"01111000110001110110111",
"01111000101001001100100",
"01111000100000100010101",
"01111000010111111001000",
"01111000001111001111111",
"01111000000110100111001",
"01110111111101111110110",
"01110111110101010110111",
"01110111101100101111010",
"01110111100100001000001",
"01110111011011100001011",
"01110111010010111011000",
"01110111001010010101000",
"01110111000001101111011",
"01110110111001001010001",
"01110110110000100101011",
"01110110101000000001000",
"01110110011111011100111",
"01110110010110111001010",
"01110110001110010110000",
"01110110000101110011010",
"01110101111101010000110",
"01110101110100101110101",
"01110101101100001101000",
"01110101100011101011110",
"01110101011011001010110",
"01110101010010101010010",
"01110101001010001010001",
"01110101000001101010011",
"01110100111001001011000",
"01110100110000101100001",
"01110100101000001101100",
"01110100011111101111010",
"01110100010111010001100",
"01110100001110110100000",
"01110100000110010111000",
"01110011111101111010011",
"01110011110101011110001",
"01110011101101000010001",
"01110011100100100110101",
"01110011011100001011100",
"01110011010011110000110",
"01110011001011010110011",
"01110011000010111100100",
"01110010111010100010111",
"01110010110010001001101",
"01110010101001110000110",
"01110010100001011000011",
"01110010011001000000010",
"01110010010000101000100",
"01110010001000010001010",
"01110001111111111010010",
"01110001110111100011101",
"01110001101111001101100",
"01110001100110110111101",
"01110001011110100010010",
"01110001010110001101001",
"01110001001101111000100",
"01110001000101100100001",
"01110000111101010000010",
"01110000110100111100101",
"01110000101100101001011",
"01110000100100010110101",
"01110000011100000100001",
"01110000010011110010001",
"01110000001011100000011",
"01110000000011001111000",
"01101111111010111110001",
"01101111110010101101100",
"01101111101010011101010",
"01101111100010001101100",
"01101111011001111110000",
"01101111010001101110111",
"01101111001001100000001",
"01101111000001010001110",
"01101110111001000011110",
"01101110110000110110001",
"01101110101000101000111",
"01101110100000011100000",
"01101110011000001111011",
"01101110010000000011010",
"01101110000111110111100",
"01101101111111101100000",
"01101101110111100001000",
"01101101101111010110010",
"01101101100111001011111",
"01101101011111000001111",
"01101101010110111000010",
"01101101001110101111001",
"01101101000110100110001",
"01101100111110011101101",
"01101100110110010101100",
"01101100101110001101110",
"01101100100110000110010",
"01101100011101111111001",
"01101100010101111000100",
"01101100001101110010001",
"01101100000101101100001",
"01101011111101100110100",
"01101011110101100001010",
"01101011101101011100010",
"01101011100101010111110",
"01101011011101010011100",
"01101011010101001111101",
"01101011001101001100010",
"01101011000101001001001",
"01101010111101000110010",
"01101010110101000011111",
"01101010101101000001111",
"01101010100101000000001",
"01101010011100111110110",
"01101010010100111101110",
"01101010001100111101001",
"01101010000100111100111",
"01101001111100111100111",
"01101001110100111101011",
"01101001101100111110001",
"01101001100100111111010",
"01101001011101000000110",
"01101001010101000010100",
"01101001001101000100110",
"01101001000101000111010",
"01101000111101001010001",
"01101000110101001101011",
"01101000101101010001000",
"01101000100101010100111",
"01101000011101011001001",
"01101000010101011101110",
"01101000001101100010110",
"01101000000101101000001",
"01100111111101101101110",
"01100111110101110011111",
"01100111101101111010001",
"01100111100110000000111",
"01100111011110001000000",
"01100111010110001111011",
"01100111001110010111001",
"01100111000110011111010",
"01100110111110100111101",
"01100110110110110000100",
"01100110101110111001101",
"01100110100111000011001",
"01100110011111001100111",
"01100110010111010111001",
"01100110001111100001101",
"01100110000111101100100",
"01100101111111110111101",
"01100101111000000011001",
"01100101110000001111000",
"01100101101000011011010",
"01100101100000100111111",
"01100101011000110100110",
"01100101010001000010000",
"01100101001001001111100",
"01100101000001011101100",
"01100100111001101011110",
"01100100110001111010011",
"01100100101010001001010",
"01100100100010011000100",
"01100100011010101000001",
"01100100010010111000001",
"01100100001011001000011",
"01100100000011011001000",
"01100011111011101010000",
"01100011110011111011010",
"01100011101100001100111",
"01100011100100011110111",
"01100011011100110001001",
"01100011010101000011110",
"01100011001101010110110",
"01100011000101101010000",
"01100010111101111101101",
"01100010110110010001101",
"01100010101110100110000",
"01100010100110111010101",
"01100010011111001111100",
"01100010010111100100111",
"01100010001111111010100",
"01100010001000010000100",
"01100010000000100110110",
"01100001111000111101011",
"01100001110001010100011",
"01100001101001101011101",
"01100001100010000011010",
"01100001011010011011001",
"01100001010010110011011",
"01100001001011001100000",
"01100001000011100101000",
"01100000111011111110010",
"01100000110100010111110",
"01100000101100110001110",
"01100000100101001100000",
"01100000011101100110100",
"01100000010110000001011",
"01100000001110011100101",
"01100000000110111000001",
"01011111111111010100000",
"01011111110111110000010",
"01011111110000001100110",
"01011111101000101001101",
"01011111100001000110110",
"01011111011001100100010",
"01011111010010000010000",
"01011111001010100000001",
"01011111000010111110101",
"01011110111011011101011",
"01011110110011111100100",
"01011110101100011011111",
"01011110100100111011101",
"01011110011101011011110",
"01011110010101111100001",
"01011110001110011100111",
"01011110000110111101111",
"01011101111111011111010",
"01011101111000000000111",
"01011101110000100010111",
"01011101101001000101001",
"01011101100001100111110",
"01011101011010001010110",
"01011101010010101110000",
"01011101001011010001101",
"01011101000011110101100",
"01011100111100011001101",
"01011100110100111110010",
"01011100101101100011000",
"01011100100110001000010",
"01011100011110101101101",
"01011100010111010011100",
"01011100001111111001100",
"01011100001000100000000",
"01011100000001000110110",
"01011011111001101101110",
"01011011110010010101001",
"01011011101010111100110",
"01011011100011100100110",
"01011011011100001101001",
"01011011010100110101110",
"01011011001101011110101",
"01011011000110000111111",
"01011010111110110001011",
"01011010110111011011010",
"01011010110000000101100",
"01011010101000101111111",
"01011010100001011010110",
"01011010011010000101111",
"01011010010010110001010",
"01011010001011011101000",
"01011010000100001001000",
"01011001111100110101011",
"01011001110101100010000",
"01011001101110001110111",
"01011001100110111100001",
"01011001011111101001110",
"01011001011000010111101",
"01011001010001000101111",
"01011001001001110100010",
"01011001000010100011001",
"01011000111011010010010",
"01011000110100000001101",
"01011000101100110001011",
"01011000100101100001011",
"01011000011110010001101",
"01011000010111000010011",
"01011000001111110011010",
"01011000001000100100100",
"01011000000001010110000",
"01010111111010000111111",
"01010111110010111010000",
"01010111101011101100100",
"01010111100100011111010",
"01010111011101010010010",
"01010111010110000101101",
"01010111001110111001010",
"01010111000111101101010",
"01010111000000100001100",
"01010110111001010110001",
"01010110110010001011000",
"01010110101011000000001",
"01010110100011110101101",
"01010110011100101011011",
"01010110010101100001011",
"01010110001110010111110",
"01010110000111001110011",
"01010110000000000101011",
"01010101111000111100101",
"01010101110001110100001",
"01010101101010101100000",
"01010101100011100100001",
"01010101011100011100101",
"01010101010101010101011",
"01010101001110001110011",
"01010101000111000111110",
"01010101000000000001011",
"01010100111000111011010",
"01010100110001110101100",
"01010100101010110000000",
"01010100100011101010111",
"01010100011100100101111",
"01010100010101100001011",
"01010100001110011101000",
"01010100000111011001000",
"01010100000000010101010",
"01010011111001010001111",
"01010011110010001110110",
"01010011101011001011111",
"01010011100100001001010",
"01010011011101000111000",
"01010011010110000101001",
"01010011001111000011011",
"01010011001000000010000",
"01010011000001000000111",
"01010010111010000000001",
"01010010110010111111101",
"01010010101011111111011",
"01010010100100111111011",
"01010010011101111111110",
"01010010010111000000011",
"01010010010000000001011",
"01010010001001000010100",
"01010010000010000100001",
"01010001111011000101111",
"01010001110100001000000",
"01010001101101001010010",
"01010001100110001101000",
"01010001011111001111111",
"01010001011000010011001",
"01010001010001010110101",
"01010001001010011010100",
"01010001000011011110100",
"01010000111100100010111",
"01010000110101100111100",
"01010000101110101100100",
"01010000100111110001110",
"01010000100000110111010",
"01010000011001111101000",
"01010000010011000011001",
"01010000001100001001100",
"01010000000101010000001",
"01001111111110010111000",
"01001111110111011110010",
"01001111110000100101110",
"01001111101001101101100",
"01001111100010110101100",
"01001111011011111101111",
"01001111010101000110100",
"01001111001110001111011",
"01001111000111011000101",
"01001111000000100010000",
"01001110111001101011110",
"01001110110010110101110",
"01001110101100000000001",
"01001110100101001010101",
"01001110011110010101100",
"01001110010111100000101",
"01001110010000101100001",
"01001110001001110111110",
"01001110000011000011110",
"01001101111100010000000",
"01001101110101011100100",
"01001101101110101001011",
"01001101100111110110011",
"01001101100001000011110",
"01001101011010010001011",
"01001101010011011111010",
"01001101001100101101100",
"01001101000101111100000",
"01001100111111001010110",
"01001100111000011001110",
"01001100110001101001000",
"01001100101010111000100",
"01001100100100001000011",
"01001100011101011000100",
"01001100010110101000111",
"01001100001111111001100",
"01001100001001001010100",
"01001100000010011011101",
"01001011111011101101001",
"01001011110100111110111",
"01001011101110010000111",
"01001011100111100011010",
"01001011100000110101110",
"01001011011010001000101",
"01001011010011011011110",
"01001011001100101111001",
"01001011000110000010110",
"01001010111111010110101",
"01001010111000101010111",
"01001010110001111111010",
"01001010101011010100000",
"01001010100100101001000",
"01001010011101111110010",
"01001010010111010011111",
"01001010010000101001101",
"01001010001001111111110",
"01001010000011010110000",
"01001001111100101100101",
"01001001110110000011100",
"01001001101111011010101",
"01001001101000110010001",
"01001001100010001001110",
"01001001011011100001110",
"01001001010100111001111",
"01001001001110010010011",
"01001001000111101011001",
"01001001000001000100001",
"01001000111010011101011",
"01001000110011110111000",
"01001000101101010000110",
"01001000100110101010111",
"01001000100000000101001",
"01001000011001011111110",
"01001000010010111010101",
"01001000001100010101110",
"01001000000101110001001",
"01000111111111001100110",
"01000111111000101000101",
"01000111110010000100111",
"01000111101011100001010",
"01000111100100111110000",
"01000111011110011011000",
"01000111010111111000001",
"01000111010001010101101",
"01000111001010110011011",
"01000111000100010001011",
"01000110111101101111110",
"01000110110111001110010",
"01000110110000101101000",
"01000110101010001100000",
"01000110100011101011011",
"01000110011101001010111",
"01000110010110101010110",
"01000110010000001010111",
"01000110001001101011010",
"01000110000011001011110",
"01000101111100101100101",
"01000101110110001101110",
"01000101101111101111001",
"01000101101001010000110",
"01000101100010110010101",
"01000101011100010100111",
"01000101010101110111010",
"01000101001111011001111",
"01000101001000111100111",
"01000101000010100000000",
"01000100111100000011011",
"01000100110101100111001",
"01000100101111001011000",
"01000100101000101111010",
"01000100100010010011110",
"01000100011011111000011",
"01000100010101011101011",
"01000100001111000010101",
"01000100001000101000000",
"01000100000010001101110",
"01000011111011110011110",
"01000011110101011010000",
"01000011101111000000100",
"01000011101000100111010",
"01000011100010001110010",
"01000011011011110101011",
"01000011010101011100111",
"01000011001111000100101",
"01000011001000101100101",
"01000011000010010100111",
"01000010111011111101011",
"01000010110101100110001",
"01000010101111001111001",
"01000010101000111000011",
"01000010100010100001111",
"01000010011100001011101",
"01000010010101110101101",
"01000010001111011111111",
"01000010001001001010011",
"01000010000010110101001",
"01000001111100100000001",
"01000001110110001011011",
"01000001101111110110111",
"01000001101001100010101",
"01000001100011001110101",
"01000001011100111010111",
"01000001010110100111011",
"01000001010000010100001",
"01000001001010000001001",
"01000001000011101110010",
"01000000111101011011110",
"01000000110111001001100",
"01000000110000110111100",
"01000000101010100101101",
"01000000100100010100001",
"01000000011110000010111",
"01000000010111110001110",
"01000000010001100001000",
"01000000001011010000011",
"01000000000101000000001",
"00111111111110110000000",
"00111111111000100000010",
"00111111110010010000101",
"00111111101100000001010",
"00111111100101110010001",
"00111111011111100011010",
"00111111011001010100110",
"00111111010011000110011",
"00111111001100111000010",
"00111111000110101010011",
"00111111000000011100101",
"00111110111010001111010",
"00111110110100000010001",
"00111110101101110101010",
"00111110100111101000100",
"00111110100001011100001",
"00111110011011001111111",
"00111110010101000100000",
"00111110001110111000010",
"00111110001000101100110",
"00111110000010100001100",
"00111101111100010110100",
"00111101110110001011110",
"00111101110000000001010",
"00111101101001110111000",
"00111101100011101101000",
"00111101011101100011001",
"00111101010111011001101",
"00111101010001010000010",
"00111101001011000111001",
"00111101000100111110011",
"00111100111110110101110",
"00111100111000101101011",
"00111100110010100101010",
"00111100101100011101011",
"00111100100110010101101",
"00111100100000001110010",
"00111100011010000111000",
"00111100010100000000001",
"00111100001101111001011",
"00111100000111110010111",
"00111100000001101100101",
"00111011111011100110101",
"00111011110101100000111",
"00111011101111011011011",
"00111011101001010110000",
"00111011100011010001000",
"00111011011101001100001",
"00111011010111000111100",
"00111011010001000011001",
"00111011001010111111000",
"00111011000100111011001",
"00111010111110110111011",
"00111010111000110100000",
"00111010110010110000110",
"00111010101100101101110",
"00111010100110101011001",
"00111010100000101000100",
"00111010011010100110010",
"00111010010100100100010",
"00111010001110100010011",
"00111010001000100000111",
"00111010000010011111100",
"00111001111100011110011",
"00111001110110011101100",
"00111001110000011100111",
"00111001101010011100011",
"00111001100100011100001",
"00111001011110011100010",
"00111001011000011100100",
"00111001010010011101000",
"00111001001100011101101",
"00111001000110011110101",
"00111001000000011111110",
"00111000111010100001010",
"00111000110100100010111",
"00111000101110100100110",
"00111000101000100110110",
"00111000100010101001001",
"00111000011100101011101",
"00111000010110101110011",
"00111000010000110001011",
"00111000001010110100101",
"00111000000100111000001",
"00110111111110111011110",
"00110111111000111111101",
"00110111110011000011110",
"00110111101101001000001",
"00110111100111001100110",
"00110111100001010001100",
"00110111011011010110101",
"00110111010101011011111",
"00110111001111100001011",
"00110111001001100111000",
"00110111000011101101000",
"00110110111101110011001",
"00110110110111111001100",
"00110110110010000000001",
"00110110101100000110111",
"00110110100110001110000",
"00110110100000010101010",
"00110110011010011100110",
"00110110010100100100100",
"00110110001110101100011",
"00110110001000110100100",
"00110110000010111101000",
"00110101111101000101100",
"00110101110111001110011",
"00110101110001010111100",
"00110101101011100000110",
"00110101100101101010010",
"00110101011111110011111",
"00110101011001111101111",
"00110101010100001000000",
"00110101001110010010011",
"00110101001000011101000",
"00110101000010100111111",
"00110100111100110010111",
"00110100110110111110001",
"00110100110001001001101",
"00110100101011010101010",
"00110100100101100001010",
"00110100011111101101011",
"00110100011001111001110",
"00110100010100000110010",
"00110100001110010011000",
"00110100001000100000000",
"00110100000010101101010",
"00110011111100111010110",
"00110011110111001000011",
"00110011110001010110010",
"00110011101011100100011",
"00110011100101110010101",
"00110011100000000001010",
"00110011011010010000000",
"00110011010100011110111",
"00110011001110101110001",
"00110011001000111101100",
"00110011000011001101001",
"00110010111101011101000",
"00110010110111101101000",
"00110010110001111101010",
"00110010101100001101110",
"00110010100110011110011",
"00110010100000101111010",
"00110010011011000000011",
"00110010010101010001110",
"00110010001111100011010",
"00110010001001110101000",
"00110010000100000111000",
"00110001111110011001010",
"00110001111000101011101",
"00110001110010111110010",
"00110001101101010001001",
"00110001100111100100001",
"00110001100001110111011",
"00110001011100001010111",
"00110001010110011110100",
"00110001010000110010011",
"00110001001011000110100",
"00110001000101011010110",
"00110000111111101111011",
"00110000111010000100001",
"00110000110100011001000",
"00110000101110101110001",
"00110000101001000011100",
"00110000100011011001001",
"00110000011101101110111",
"00110000011000000100111",
"00110000010010011011001",
"00110000001100110001100",
"00110000000111001000001",
"00110000000001011111000",
"00101111111011110110001",
"00101111110110001101011",
"00101111110000100100110",
"00101111101010111100100",
"00101111100101010100011",
"00101111011111101100100",
"00101111011010000100110",
"00101111010100011101010",
"00101111001110110110000",
"00101111001001001110111",
"00101111000011101000000",
"00101110111110000001011",
"00101110111000011010111",
"00101110110010110100101",
"00101110101101001110101",
"00101110100111101000111",
"00101110100010000011001",
"00101110011100011101110",
"00101110010110111000100",
"00101110010001010011100",
"00101110001011101110110",
"00101110000110001010001",
"00101110000000100101110",
"00101101111011000001101",
"00101101110101011101101",
"00101101101111111001111",
"00101101101010010110010",
"00101101100100110010111",
"00101101011111001111110",
"00101101011001101100110",
"00101101010100001010000",
"00101101001110100111100",
"00101101001001000101001",
"00101101000011100011000",
"00101100111110000001000",
"00101100111000011111010",
"00101100110010111101110",
"00101100101101011100100",
"00101100100111111011011",
"00101100100010011010011",
"00101100011100111001101",
"00101100010111011001001",
"00101100010001111000111",
"00101100001100011000110",
"00101100000110111000110",
"00101100000001011001001",
"00101011111011111001101",
"00101011110110011010010",
"00101011110000111011001",
"00101011101011011100010",
"00101011100101111101100",
"00101011100000011111000",
"00101011011011000000110",
"00101011010101100010101",
"00101011010000000100101",
"00101011001010100111000",
"00101011000101001001100",
"00101010111111101100001",
"00101010111010001111000",
"00101010110100110010001",
"00101010101111010101011",
"00101010101001111000111",
"00101010100100011100101",
"00101010011111000000100",
"00101010011001100100100",
"00101010010100001000111",
"00101010001110101101010",
"00101010001001010010000",
"00101010000011110110111",
"00101001111110011011111",
"00101001111001000001001",
"00101001110011100110101",
"00101001101110001100010",
"00101001101000110010001",
"00101001100011011000010",
"00101001011101111110100",
"00101001011000100100111",
"00101001010011001011100",
"00101001001101110010011",
"00101001001000011001011",
"00101001000011000000101",
"00101000111101101000000",
"00101000111000001111101",
"00101000110010110111100",
"00101000101101011111100",
"00101000101000000111101",
"00101000100010110000001",
"00101000011101011000101",
"00101000011000000001100",
"00101000010010101010011",
"00101000001101010011101",
"00101000000111111101000",
"00101000000010100110100",
"00100111111101010000010",
"00100111110111111010010",
"00100111110010100100011",
"00100111101101001110110",
"00100111100111111001010",
"00100111100010100100000",
"00100111011101001110111",
"00100111010111111010000",
"00100111010010100101010",
"00100111001101010000110",
"00100111000111111100011",
"00100111000010101000010",
"00100110111101010100011",
"00100110111000000000101",
"00100110110010101101000",
"00100110101101011001101",
"00100110101000000110100",
"00100110100010110011100",
"00100110011101100000110",
"00100110011000001110001",
"00100110010010111011101",
"00100110001101101001100",
"00100110001000010111011",
"00100110000011000101101",
"00100101111101110011111",
"00100101111000100010100",
"00100101110011010001001",
"00100101101110000000001",
"00100101101000101111001",
"00100101100011011110100",
"00100101011110001110000",
"00100101011000111101101",
"00100101010011101101100",
"00100101001110011101100",
"00100101001001001101110",
"00100101000011111110001",
"00100100111110101110110",
"00100100111001011111100",
"00100100110100010000100",
"00100100101111000001110",
"00100100101001110011000",
"00100100100100100100101",
"00100100011111010110010",
"00100100011010001000010",
"00100100010100111010011",
"00100100001111101100101",
"00100100001010011111001",
"00100100000101010001110",
"00100100000000000100101",
"00100011111010110111101",
"00100011110101101010110",
"00100011110000011110010",
"00100011101011010001110",
"00100011100110000101100",
"00100011100000111001100",
"00100011011011101101101",
"00100011010110100010000",
"00100011010001010110100",
"00100011001100001011001",
"00100011000111000000000",
"00100011000001110101001",
"00100010111100101010011",
"00100010110111011111110",
"00100010110010010101011",
"00100010101101001011001",
"00100010101000000001001",
"00100010100010110111010",
"00100010011101101101101",
"00100010011000100100001",
"00100010010011011010111",
"00100010001110010001110",
"00100010001001001000111",
"00100010000100000000001",
"00100001111110110111100",
"00100001111001101111001",
"00100001110100100110111",
"00100001101111011110111",
"00100001101010010111000",
"00100001100101001111011",
"00100001100000000111111",
"00100001011011000000101",
"00100001010101111001100",
"00100001010000110010101",
"00100001001011101011111",
"00100001000110100101010",
"00100001000001011110111",
"00100000111100011000101",
"00100000110111010010101",
"00100000110010001100110",
"00100000101101000111000",
"00100000101000000001100",
"00100000100010111100010",
"00100000011101110111001",
"00100000011000110010001",
"00100000010011101101011",
"00100000001110101000110",
"00100000001001100100011",
"00100000000100100000001",
"00011111111111011100000",
"00011111111010011000001",
"00011111110101010100011",
"00011111110000010000111",
"00011111101011001101100",
"00011111100110001010011",
"00011111100001000111011",
"00011111011100000100100",
"00011111010111000001111",
"00011111010001111111011",
"00011111001100111101001",
"00011111000111111011000",
"00011111000010111001000",
"00011110111101110111010",
"00011110111000110101101",
"00011110110011110100010",
"00011110101110110011000",
"00011110101001110010000",
"00011110100100110001000",
"00011110011111110000011",
"00011110011010101111110",
"00011110010101101111100",
"00011110010000101111010",
"00011110001011101111010",
"00011110000110101111011",
"00011110000001101111110",
"00011101111100110000010",
"00011101110111110000111",
"00011101110010110001110",
"00011101101101110010111",
"00011101101000110100000",
"00011101100011110101011",
"00011101011110110111000",
"00011101011001111000110",
"00011101010100111010101",
"00011101001111111100101",
"00011101001010111110111",
"00011101000110000001011",
"00011101000001000011111",
"00011100111100000110101",
"00011100110111001001101",
"00011100110010001100110",
"00011100101101010000000",
"00011100101000010011100",
"00011100100011010111001",
"00011100011110011010111",
"00011100011001011110111",
"00011100010100100011000",
"00011100001111100111010",
"00011100001010101011110",
"00011100000101110000011",
"00011100000000110101010",
"00011011111011111010010",
"00011011110110111111011",
"00011011110010000100110",
"00011011101101001010010",
"00011011101000001111111",
"00011011100011010101110",
"00011011011110011011110",
"00011011011001100010000",
"00011011010100101000011",
"00011011001111101110111",
"00011011001010110101100",
"00011011000101111100011",
"00011011000001000011100",
"00011010111100001010101",
"00011010110111010010000",
"00011010110010011001100",
"00011010101101100001010",
"00011010101000101001001",
"00011010100011110001001",
"00011010011110111001011",
"00011010011010000001110",
"00011010010101001010010",
"00011010010000010011000",
"00011010001011011011111",
"00011010000110100101000",
"00011010000001101110001",
"00011001111100110111100",
"00011001111000000001001",
"00011001110011001010111",
"00011001101110010100110",
"00011001101001011110110",
"00011001100100101001000",
"00011001011111110011011",
"00011001011010111101111",
"00011001010110001000101",
"00011001010001010011100",
"00011001001100011110100",
"00011001000111101001110",
"00011001000010110101001",
"00011000111110000000110",
"00011000111001001100011",
"00011000110100011000010",
"00011000101111100100011",
"00011000101010110000100",
"00011000100101111100111",
"00011000100001001001011",
"00011000011100010110001",
"00011000010111100011000",
"00011000010010110000000",
"00011000001101111101010",
"00011000001001001010100",
"00011000000100011000001",
"00010111111111100101110",
"00010111111010110011101",
"00010111110110000001101",
"00010111110001001111110",
"00010111101100011110001",
"00010111100111101100101",
"00010111100010111011010",
"00010111011110001010001",
"00010111011001011001001",
"00010111010100101000010",
"00010111001111110111100",
"00010111001011000111000",
"00010111000110010110101",
"00010111000001100110100",
"00010110111100110110011",
"00010110111000000110100",
"00010110110011010110111",
"00010110101110100111010",
"00010110101001110111111",
"00010110100101001000101",
"00010110100000011001101",
"00010110011011101010101",
"00010110010110111011111",
"00010110010010001101011",
"00010110001101011110111",
"00010110001000110000101",
"00010110000100000010100",
"00010101111111010100101",
"00010101111010100110110",
"00010101110101111001001",
"00010101110001001011101",
"00010101101100011110011",
"00010101100111110001010",
"00010101100011000100010",
"00010101011110010111011",
"00010101011001101010110",
"00010101010100111110010",
"00010101010000010001111",
"00010101001011100101101",
"00010101000110111001101",
"00010101000010001101110",
"00010100111101100010000",
"00010100111000110110100",
"00010100110100001011001",
"00010100101111011111111",
"00010100101010110100110",
"00010100100110001001111",
"00010100100001011111000",
"00010100011100110100100",
"00010100011000001010000",
"00010100010011011111110",
"00010100001110110101100",
"00010100001010001011101",
"00010100000101100001110",
"00010100000000111000001",
"00010011111100001110100",
"00010011110111100101010",
"00010011110010111100000",
"00010011101110010011000",
"00010011101001101010001",
"00010011100101000001011",
"00010011100000011000110",
"00010011011011110000011",
"00010011010111001000001",
"00010011010010100000000",
"00010011001101111000000",
"00010011001001010000010",
"00010011000100101000101",
"00010011000000000001001",
"00010010111011011001110",
"00010010110110110010101",
"00010010110010001011100",
"00010010101101100100101",
"00010010101000111110000",
"00010010100100010111011",
"00010010011111110001000",
"00010010011011001010110",
"00010010010110100100101",
"00010010010001111110110",
"00010010001101011000111",
"00010010001000110011010",
"00010010000100001101110",
"00010001111111101000100",
"00010001111011000011010",
"00010001110110011110010",
"00010001110001111001011",
"00010001101101010100101",
"00010001101000110000001",
"00010001100100001011110",
"00010001011111100111011",
"00010001011011000011011",
"00010001010110011111011",
"00010001010001111011101",
"00010001001101010111111",
"00010001001000110100011",
"00010001000100010001001",
"00010000111111101101111",
"00010000111011001010111",
"00010000110110101000000",
"00010000110010000101010",
"00010000101101100010101",
"00010000101001000000001",
"00010000100100011101111",
"00010000011111111011110",
"00010000011011011001110",
"00010000010110110111111",
"00010000010010010110010",
"00010000001101110100110",
"00010000001001010011011",
"00010000000100110010001",
"00010000000000010001000",
"00001111111011110000001",
"00001111110111001111010",
"00001111110010101110101",
"00001111101110001110001",
"00001111101001101101111",
"00001111100101001101101",
"00001111100000101101101",
"00001111011100001101110",
"00001111010111101110000",
"00001111010011001110011",
"00001111001110101111000",
"00001111001010001111101",
"00001111000101110000100",
"00001111000001010001100",
"00001110111100110010101",
"00001110111000010100000",
"00001110110011110101011",
"00001110101111010111000",
"00001110101010111000110",
"00001110100110011010101",
"00001110100001111100110",
"00001110011101011110111",
"00001110011001000001010",
"00001110010100100011110",
"00001110010000000110011",
"00001110001011101001001",
"00001110000111001100000",
"00001110000010101111001",
"00001101111110010010011",
"00001101111001110101110",
"00001101110101011001010",
"00001101110000111100111",
"00001101101100100000101",
"00001101101000000100101",
"00001101100011101000110",
"00001101011111001101000",
"00001101011010110001011",
"00001101010110010101111",
"00001101010001111010100",
"00001101001101011111011",
"00001101001001000100011",
"00001101000100101001100",
"00001101000000001110110",
"00001100111011110100001",
"00001100110111011001101",
"00001100110010111111011",
"00001100101110100101010",
"00001100101010001011001",
"00001100100101110001011",
"00001100100001010111101",
"00001100011100111110000",
"00001100011000100100101",
"00001100010100001011010",
"00001100001111110010001",
"00001100001011011001001",
"00001100000111000000010",
"00001100000010100111100",
"00001011111110001111000",
"00001011111001110110100",
"00001011110101011110010",
"00001011110001000110001",
"00001011101100101110001",
"00001011101000010110010",
"00001011100011111110100",
"00001011011111100110111",
"00001011011011001111100",
"00001011010110111000010",
"00001011010010100001000",
"00001011001110001010000",
"00001011001001110011001",
"00001011000101011100100",
"00001011000001000101111",
"00001010111100101111100",
"00001010111000011001001",
"00001010110100000011000",
"00001010101111101101000",
"00001010101011010111001",
"00001010100111000001011",
"00001010100010101011110",
"00001010011110010110011",
"00001010011010000001000",
"00001010010101101011111",
"00001010010001010110111",
"00001010001101000010000",
"00001010001000101101010",
"00001010000100011000101",
"00001010000000000100001",
"00001001111011101111111",
"00001001110111011011101",
"00001001110011000111101",
"00001001101110110011110",
"00001001101010100000000",
"00001001100110001100011",
"00001001100001111000111",
"00001001011101100101100",
"00001001011001010010010",
"00001001010100111111010",
"00001001010000101100010",
"00001001001100011001100",
"00001001001000000110111",
"00001001000011110100011",
"00001000111111100010000",
"00001000111011001111110",
"00001000110110111101101",
"00001000110010101011110",
"00001000101110011001111",
"00001000101010001000010",
"00001000100101110110101",
"00001000100001100101010",
"00001000011101010100000",
"00001000011001000010111",
"00001000010100110001111",
"00001000010000100001000",
"00001000001100010000011",
"00001000000111111111110",
"00001000000011101111010",
"00000111111111011111000",
"00000111111011001110111",
"00000111110110111110110",
"00000111110010101110111",
"00000111101110011111001",
"00000111101010001111100",
"00000111100110000000001",
"00000111100001110000110",
"00000111011101100001100",
"00000111011001010010100",
"00000111010101000011100",
"00000111010000110100110",
"00000111001100100110000",
"00000111001000010111100",
"00000111000100001001001",
"00000110111111111010111",
"00000110111011101100110",
"00000110110111011110110",
"00000110110011010000111",
"00000110101111000011010",
"00000110101010110101101",
"00000110100110101000001",
"00000110100010011010111",
"00000110011110001101101",
"00000110011010000000101",
"00000110010101110011110",
"00000110010001100111000",
"00000110001101011010011",
"00000110001001001101111",
"00000110000101000001100",
"00000110000000110101010",
"00000101111100101001001",
"00000101111000011101001",
"00000101110100010001011",
"00000101110000000101101",
"00000101101011111010000",
"00000101100111101110101",
"00000101100011100011011",
"00000101011111011000001",
"00000101011011001101001",
"00000101010111000010010",
"00000101010010110111100",
"00000101001110101100111",
"00000101001010100010011",
"00000101000110011000000",
"00000101000010001101110",
"00000100111110000011101",
"00000100111001111001101",
"00000100110101101111111",
"00000100110001100110001",
"00000100101101011100100",
"00000100101001010011001",
"00000100100101001001110",
"00000100100001000000101",
"00000100011100110111101",
"00000100011000101110101",
"00000100010100100101111",
"00000100010000011101010",
"00000100001100010100110",
"00000100001000001100011",
"00000100000100000100001",
"00000011111111111100000",
"00000011111011110100000",
"00000011110111101100001",
"00000011110011100100011",
"00000011101111011100110",
"00000011101011010101010",
"00000011100111001101111",
"00000011100011000110110",
"00000011011110111111101",
"00000011011010111000101",
"00000011010110110001111",
"00000011010010101011001",
"00000011001110100100101",
"00000011001010011110001",
"00000011000110010111111",
"00000011000010010001110",
"00000010111110001011101",
"00000010111010000101110",
"00000010110110000000000",
"00000010110001111010011",
"00000010101101110100110",
"00000010101001101111011",
"00000010100101101010001",
"00000010100001100101000",
"00000010011101100000000",
"00000010011001011011001",
"00000010010101010110011",
"00000010010001010001110",
"00000010001101001101010",
"00000010001001001000111",
"00000010000101000100101",
"00000010000001000000100",
"00000001111100111100100",
"00000001111000111000101",
"00000001110100110101000",
"00000001110000110001011",
"00000001101100101101111",
"00000001101000101010100",
"00000001100100100111010",
"00000001100000100100010",
"00000001011100100001010",
"00000001011000011110011",
"00000001010100011011110",
"00000001010000011001001",
"00000001001100010110101",
"00000001001000010100011",
"00000001000100010010001",
"00000001000000010000001",
"00000000111100001110001",
"00000000111000001100010",
"00000000110100001010101",
"00000000110000001001000",
"00000000101100000111101",
"00000000101000000110010",
"00000000100100000101001",
"00000000100000000100000",
"00000000011100000011001",
"00000000011000000010010",
"00000000010100000001101",
"00000000010000000001000",
"00000000001100000000101",
"00000000001000000000010",
"00000000000100000000001");
  constant rom2 : rom_t :=("11111111111111111111110",
"11111111100000000001100",
"11111111000000000110000",
"11111110100000001101100",
"11111110000000011000000",
"11111101100000100101100",
"11111101000000110101111",
"11111100100001001001011",
"11111100000001011111110",
"11111011100001111000111",
"11111011000010010101010",
"11111010100010110100011",
"11111010000011010110011",
"11111001100011111011011",
"11111001000100100011011",
"11111000100101001110011",
"11111000000101111100010",
"11110111100110101100111",
"11110111000111100000100",
"11110110101000010111000",
"11110110001001010000011",
"11110101101010001100110",
"11110101001011001011111",
"11110100101100001101111",
"11110100001101010010111",
"11110011101110011010100",
"11110011001111100101011",
"11110010110000110010111",
"11110010010010000011000",
"11110001110011010110011",
"11110001010100101100011",
"11110000110110000101000",
"11110000010111100000101",
"11101111111000111111001",
"11101111011010100000100",
"11101110111100000100101",
"11101110011101101011100",
"11101101111111010101001",
"11101101100001000001101",
"11101101000010110001001",
"11101100100100100011001",
"11101100000110011000001",
"11101011101000001111101",
"11101011001010001001111",
"11101010101100000111010",
"11101010001110000110111",
"11101001110000001001110",
"11101001010010001111000",
"11101000110100010111001",
"11101000010110100010000",
"11100111111000101111101",
"11100111011011000000001",
"11100110111101010011001",
"11100110011111101000110",
"11100110000010000001010",
"11100101100100011100011",
"11100101000110111010011",
"11100100101001011011000",
"11100100001011111110001",
"11100011101110100100001",
"11100011010001001100110",
"11100010110011110111111",
"11100010010110100110000",
"11100001111001010110100",
"11100001011100001001110",
"11100000111110111111110",
"11100000100001111000001",
"11100000000100110011100",
"11011111100111110001010",
"11011111001010110001111",
"11011110101101110101000",
"11011110010000111010101",
"11011101110100000010111",
"11011101010111001110000",
"11011100111010011011101",
"11011100011101101011110",
"11011100000000111110100",
"11011011100100010011110",
"11011011000111101011111",
"11011010101011000110010",
"11011010001110100011011",
"11011001110010000011001",
"11011001010101100101011",
"11011000111001001010001",
"11011000011100110001100",
"11011000000000011011101",
"11010111100100001000000",
"11010111000111110111001",
"11010110101011101000100",
"11010110001111011100110",
"11010101110011010011100",
"11010101010111001100100",
"11010100111011001000010",
"11010100011111000110100",
"11010100000011000111000",
"11010011100111001010010",
"11010011001011010000001",
"11010010101111011000011",
"11010010010011100010111",
"11010001110111110000010",
"11010001011011111111110",
"11010001000000010010001",
"11010000100100100110101",
"11010000001000111101101",
"11001111101101010111011",
"11001111010001110011011",
"11001110110110010001111",
"11001110011010110010111",
"11001101111111010110001",
"11001101100011111100000",
"11001101001000100100010",
"11001100101101001111001",
"11001100010001111100001",
"11001011110110101011110",
"11001011011011011101100",
"11001011000000010010000",
"11001010100101001000110",
"11001010001010000010000",
"11001001101110111101101",
"11001001010011111011110",
"11001000111000111100000",
"11001000011101111110110",
"11001000000011000100000",
"11000111101000001011101",
"11000111001101010101100",
"11000110110010100001110",
"11000110010111110000100",
"11000101111101000001100",
"11000101100010010100111",
"11000101000111101010101",
"11000100101101000010111",
"11000100010010011101010",
"11000011110111111001111",
"11000011011101011001001",
"11000011000010111010101",
"11000010101000011110010",
"11000010001110000100011",
"11000001110011101100111",
"11000001011001010111110",
"11000000111111000100100",
"11000000100100110100000",
"11000000001010100101101",
"10111111110000011001110",
"10111111010110001111111",
"10111110111100001000100",
"10111110100010000011010",
"10111110001000000000100",
"10111101101101111111110",
"10111101010100000001100",
"10111100111010000101011",
"10111100100000001011011",
"10111100000110010100000",
"10111011101100011110101",
"10111011010010101011100",
"10111010111000111010111",
"10111010011111001100011",
"10111010000101100000000",
"10111001101011110101111",
"10111001010010001110000",
"10111000111000101000100",
"10111000011111000101001",
"10111000000101100100001",
"10110111101100000101000",
"10110111010010101000100",
"10110110111001001101111",
"10110110011111110101100",
"10110110000110011111011",
"10110101101101001011100",
"10110101010011111001111",
"10110100111010101010010",
"10110100100001011100111",
"10110100001000010001110",
"10110011101111001000110",
"10110011010110000001110",
"10110010111100111101010",
"10110010100011111010110",
"10110010001010111010011",
"10110001110001111100001",
"10110001011001000000010",
"10110001000000000110011",
"10110000100111001110101",
"10110000001110011001000",
"10101111110101100101101",
"10101111011100110100011",
"10101111000100000101000",
"10101110101011011000010",
"10101110010010101101010",
"10101101111010000100011",
"10101101100001011101110",
"10101101001000111001000",
"10101100110000010110100",
"10101100010111110110010",
"10101011111111010111111",
"10101011100110111011111",
"10101011001110100001110",
"10101010110110001001101",
"10101010011101110011111",
"10101010000101011111111",
"10101001101101001110010",
"10101001010100111110101",
"10101000111100110001001",
"10101000100100100101011",
"10101000001100011011111",
"10100111110100010100100",
"10100111011100001111001",
"10100111000100001011111",
"10100110101100001010101",
"10100110010100001011011",
"10100101111100001110010",
"10100101100100010011001",
"10100101001100011010000",
"10100100110100100011000",
"10100100011100101101110",
"10100100000100111010110",
"10100011101101001001111",
"10100011010101011010111",
"10100010111101101101110",
"10100010100110000011000",
"10100010001110011001111",
"10100001110110110011001",
"10100001011111001110000",
"10100001000111101011000",
"10100000110000001010001",
"10100000011000101011001",
"10100000000001001110001",
"10011111101001110011000",
"10011111010010011010001",
"10011110111011000010111",
"10011110100011101101110",
"10011110001100011010101",
"10011101110101001001100",
"10011101011101111010011",
"10011101000110101101000",
"10011100101111100001110",
"10011100011000011000011",
"10011100000001010001000",
"10011011101010001011101",
"10011011010011001000000",
"10011010111100000110011",
"10011010100101000110110",
"10011010001110001001001",
"10011001110111001101010",
"10011001100000010011011",
"10011001001001011011100",
"10011000110010100101011",
"10011000011011110001001",
"10011000000100111111000",
"10010111101110001110110",
"10010111010111100000010",
"10010111000000110011110",
"10010110101010001001010",
"10010110010011100000011",
"10010101111100111001101",
"10010101100110010100110",
"10010101001111110001101",
"10010100111001010000011",
"10010100100010110001000",
"10010100001100010011100",
"10010011110101111000000",
"10010011011111011110010",
"10010011001001000110011",
"10010010110010110000100",
"10010010011100011100011",
"10010010000110001010010",
"10010001101111111001110",
"10010001011001101011010",
"10010001000011011110011",
"10010000101101010011100",
"10010000010111001010011",
"10010000000001000011001",
"10001111101010111101111",
"10001111010100111010011",
"10001110111110111000100",
"10001110101000111000101",
"10001110010010111010101",
"10001101111100111110010",
"10001101100111000100000",
"10001101010001001011001",
"10001100111011010100011",
"10001100100101011111011",
"10001100001111101100000",
"10001011111001111010101",
"10001011100100001010111",
"10001011001110011101001",
"10001010111000110001000",
"10001010100011000110101",
"10001010001101011110001",
"10001001110111110111100",
"10001001100010010010011",
"10001001001100101111011",
"10001000110111001101111",
"10001000100001101110010",
"10001000001100010000011",
"10000111110110110100010",
"10000111100001011001111",
"10000111001100000001010",
"10000110110110101010011",
"10000110100001010101011",
"10000110001100000001111",
"10000101110110110000011",
"10000101100001100000100",
"10000101001100010010010",
"10000100110111000101111",
"10000100100001111011010",
"10000100001100110010010",
"10000011110111101010111",
"10000011100010100101100",
"10000011001101100001101",
"10000010111000011111100",
"10000010100011011111010",
"10000010001110100000100",
"10000001111001100011100",
"10000001100100101000100",
"10000001001111101110110",
"10000000111010110111000",
"10000000100110000000111",
"10000000010001001100011",
"01111111111100011001101",
"01111111100111101000011",
"01111111010010111001001",
"01111110111110001011011",
"01111110101001011111011",
"01111110010100110101000",
"01111110000000001100011",
"01111101101011100101010",
"01111101010111000000000",
"01111101000010011100011",
"01111100101101111010011",
"01111100011001011001111",
"01111100000100111011001",
"01111011110000011110000",
"01111011011100000010110",
"01111011000111101000111",
"01111010110011010000111",
"01111010011110111010100",
"01111010001010100101011",
"01111001110110010010010",
"01111001100010000000110",
"01111001001101110000110",
"01111000111001100010100",
"01111000100101010110000",
"01111000010001001010111",
"01110111111101000001011",
"01110111101000111001100",
"01110111010100110011010",
"01110111000000101110110",
"01110110101100101011110",
"01110110011000101010011",
"01110110000100101010110",
"01110101110000101100100",
"01110101011100101111111",
"01110101001000110101000",
"01110100110100111011100",
"01110100100001000011110",
"01110100001101001101100",
"01110011111001011001000",
"01110011100101100110000",
"01110011010001110100100",
"01110010111110000100101",
"01110010101010010110011",
"01110010010110101001101",
"01110010000010111110010",
"01110001101111010100110",
"01110001011011101100111",
"01110001001000000110010",
"01110000110100100001100",
"01110000100000111110001",
"01110000001101011100010",
"01101111111001111100000",
"01101111100110011101010",
"01101111010011000000001",
"01101110111111100100101",
"01101110101100001010100",
"01101110011000110010001",
"01101110000101011011000",
"01101101110010000101101",
"01101101011110110001101",
"01101101001011011111011",
"01101100111000001110011",
"01101100100100111111001",
"01101100010001110001010",
"01101011111110100101000",
"01101011101011011010001",
"01101011011000010000111",
"01101011000101001001001",
"01101010110010000010110",
"01101010011110111110001",
"01101010001011111010111",
"01101001111000111001001",
"01101001100101111000110",
"01101001010010111010001",
"01101000111111111100111",
"01101000101101000001000",
"01101000011010000110110",
"01101000000111001110000",
"01100111110100010110110",
"01100111100001100000111",
"01100111001110101100101",
"01100110111011111001110",
"01100110101001001000011",
"01100110010110011000011",
"01100110000011101010000",
"01100101110000111100111",
"01100101011110010001011",
"01100101001011100111011",
"01100100111000111110111",
"01100100100110010111110",
"01100100010011110001111",
"01100100000001001101111",
"01100011101110101011000",
"01100011011100001001101",
"01100011001001101001111",
"01100010110111001011011",
"01100010100100101110010",
"01100010010010010010110",
"01100001111111111000101",
"01100001101101011111111",
"01100001011011001000101",
"01100001001000110010111",
"01100000110110011110100",
"01100000100100001011101",
"01100000010001111010000",
"01011111111111101001111",
"01011111101101011011001",
"01011111011011001101111",
"01011111001001000001111",
"01011110110110110111011",
"01011110100100101110011",
"01011110010010100110110",
"01011110000000100000100",
"01011101101110011011101",
"01011101011100011000000",
"01011101001010010110001",
"01011100111000010101011",
"01011100100110010110001",
"01011100010100011000010",
"01011100000010011011110",
"01011011110000100000110",
"01011011011110100111000",
"01011011001100101110110",
"01011010111010110111110",
"01011010101001000010000",
"01011010010111001101111",
"01011010000101011011000",
"01011001110011101001100",
"01011001100001111001100",
"01011001010000001010101",
"01011000111110011101100",
"01011000101100110001011",
"01011000011011000110110",
"01011000001001011101100",
"01010111110111110101100",
"01010111100110001111000",
"01010111010100101001101",
"01010111000011000101110",
"01010110110001100011011",
"01010110100000000010010",
"01010110001110100010011",
"01010101111101000011110",
"01010101101011100110101",
"01010101011010001010110",
"01010101001000110000010",
"01010100110111010111001",
"01010100100101111111010",
"01010100010100101000110",
"01010100000011010011101",
"01010011110001111111101",
"01010011100000101101010",
"01010011001111011100000",
"01010010111110001100000",
"01010010101100111101100",
"01010010011011110000010",
"01010010001010100100010",
"01010001111001011001110",
"01010001101000010000010",
"01010001010111001000011",
"01010001000110000001101",
"01010000110100111100000",
"01010000100011110111111",
"01010000010010110101010",
"01010000000001110011101",
"01001111110000110011011",
"01001111011111110100100",
"01001111001110110110110",
"01001110111101111010010",
"01001110101100111111010",
"01001110011100000101011",
"01001110001011001100111",
"01001101111010010101100",
"01001101101001011111101",
"01001101011000101010110",
"01001101000111110111011",
"01001100110111000101001",
"01001100100110010100011",
"01001100010101100100101",
"01001100000100110110010",
"01001011110100001001010",
"01001011100011011101011",
"01001011010010110010110",
"01001011000010001001010",
"01001010110001100001010",
"01001010100000111010100",
"01001010010000010101000",
"01001001111111110000011",
"01001001101111001101100",
"01001001011110101011101",
"01001001001110001010111",
"01001000111101101011101",
"01001000101101001101011",
"01001000011100110000101",
"01001000001100010101000",
"01000111111011111010100",
"01000111101011100001011",
"01000111011011001001011",
"01000111001010110010110",
"01000110111010011101001",
"01000110101010001000110",
"01000110011001110101111",
"01000110001001100011111",
"01000101111001010011010",
"01000101101001000100000",
"01000101011000110101101",
"01000101001000101000101",
"01000100111000011100111",
"01000100101000010010011",
"01000100011000001001000",
"01000100001000000000111",
"01000011110111111001111",
"01000011100111110100001",
"01000011010111101111100",
"01000011000111101100001",
"01000010110111101010000",
"01000010100111101001000",
"01000010010111101001001",
"01000010000111101010110",
"01000001110111101101011",
"01000001100111110001001",
"01000001010111110110000",
"01000001000111111100010",
"01000000111000000011100",
"01000000101000001100000",
"01000000011000010101110",
"01000000001000100000101",
"00111111111000101100100",
"00111111101000111001110",
"00111111011001001000001",
"00111111001001010111110",
"00111110111001101000010",
"00111110101001111010010",
"00111110011010001101001",
"00111110001010100001100",
"00111101111010110110110",
"00111101101011001101010",
"00111101011011100100111",
"00111101001011111101101",
"00111100111100010111101",
"00111100101100110010110",
"00111100011101001111000",
"00111100001101101100100",
"00111011111110001011000",
"00111011101110101010110",
"00111011011111001011100",
"00111011001111101101100",
"00111011000000010000101",
"00111010110000110100111",
"00111010100001011010010",
"00111010010010000000110",
"00111010000010101000100",
"00111001110011010001001",
"00111001100011111011000",
"00111001010100100110001",
"00111001000101010010010",
"00111000110101111111011",
"00111000100110101101111",
"00111000010111011101011",
"00111000001000001110000",
"00110111111000111111110",
"00110111101001110010100",
"00110111011010100110100",
"00110111001011011011101",
"00110110111100010001110",
"00110110101101001001000",
"00110110011110000001100",
"00110110001110111011000",
"00110101111111110101100",
"00110101110000110001010",
"00110101100001101110001",
"00110101010010101011111",
"00110101000011101010111",
"00110100110100101010111",
"00110100100101101100001",
"00110100010110101110100",
"00110100000111110001110",
"00110011111000110110010",
"00110011101001111011101",
"00110011011011000010011",
"00110011001100001010000",
"00110010111101010010111",
"00110010101110011100100",
"00110010011111100111011",
"00110010010000110011011",
"00110010000010000000101",
"00110001110011001110101",
"00110001100100011101111",
"00110001010101101110001",
"00110001000110111111011",
"00110000111000010010000",
"00110000101001100101011",
"00110000011010111010000",
"00110000001100001111100",
"00101111111101100110010",
"00101111101110111101111",
"00101111100000010110101",
"00101111010001110000100",
"00101111000011001011010",
"00101110110100100111010",
"00101110100110000100010",
"00101110010111100010010",
"00101110001001000001010",
"00101101111010100001100",
"00101101101100000010101",
"00101101011101100100111",
"00101101001111001000000",
"00101101000000101100010",
"00101100110010010001101",
"00101100100011111000000",
"00101100010101011111011",
"00101100000111000111110",
"00101011111000110001001",
"00101011101010011011110",
"00101011011100000111010",
"00101011001101110011110",
"00101010111111100001010",
"00101010110001001111111",
"00101010100010111111100",
"00101010010100110000001",
"00101010000110100001101",
"00101001111000010100010",
"00101001101010001000000",
"00101001011011111100101",
"00101001001101110010011",
"00101000111111101001000",
"00101000110001100000110",
"00101000100011011001101",
"00101000010101010011011",
"00101000000111001110000",
"00100111111001001001110",
"00100111101011000110011",
"00100111011101000100001",
"00100111001111000011000",
"00100111000001000010110",
"00100110110011000011011",
"00100110100101000101001",
"00100110010111001000000",
"00100110001001001011101",
"00100101111011010000010",
"00100101101101010110000",
"00100101011111011100101",
"00100101010001100100010",
"00100101000011101101000",
"00100100110101110110110",
"00100100101000000001010",
"00100100011010001100111",
"00100100001100011001100",
"00100011111110100110111",
"00100011110000110101011",
"00100011100011000101000",
"00100011010101010101100",
"00100011000111100110111",
"00100010111001111001010",
"00100010101100001100101",
"00100010011110100001000",
"00100010010000110110011",
"00100010000011001100110",
"00100001110101100011110",
"00100001100111111100001",
"00100001011010010101001",
"00100001001100101111011",
"00100000111111001010011",
"00100000110001100110100",
"00100000100100000011011",
"00100000010110100001011",
"00100000001001000000010",
"00011111111011100000000",
"00011111101110000000111",
"00011111100000100010100",
"00011111010011000101011",
"00011111000101101001000",
"00011110111000001101100",
"00011110101010110011001",
"00011110011101011001100",
"00011110010000000000111",
"00011110000010101001010",
"00011101110101010010100",
"00011101100111111100101",
"00011101011010100111111",
"00011101001101010011111",
"00011101000000000000111",
"00011100110010101110111",
"00011100100101011101110",
"00011100011000001101011",
"00011100001010111110010",
"00011011111101101111111",
"00011011110000100010011",
"00011011100011010101110",
"00011011010110001010010",
"00011011001000111111100",
"00011010111011110101111",
"00011010101110101100111",
"00011010100001100100111",
"00011010010100011101111",
"00011010000111010111111",
"00011001111010010010101",
"00011001101101001110011",
"00011001100000001011000",
"00011001010011001000100",
"00011001000110000111000",
"00011000111001000110011",
"00011000101100000110100",
"00011000011111000111110",
"00011000010010001001110",
"00011000000101001100110",
"00010111111000010000100",
"00010111101011010101001",
"00010111011110011010110",
"00010111010001100001010",
"00010111000100101000101",
"00010110110111110001001",
"00010110101010111010011",
"00010110011110000100010",
"00010110010001001111011",
"00010110000100011011010",
"00010101110111100111111",
"00010101101010110101100",
"00010101011110000100001",
"00010101010001010011100",
"00010101000100100011101",
"00010100110111110100111",
"00010100101011000110111",
"00010100011110011001110",
"00010100010001101101100",
"00010100000101000010001",
"00010011111000010111111",
"00010011101011101110001",
"00010011011111000101100",
"00010011010010011101101",
"00010011000101110110101",
"00010010111001010000100",
"00010010101100101011001",
"00010010100000000110101",
"00010010010011100011010",
"00010010000111000000101",
"00010001111010011110101",
"00010001101101111101101",
"00010001100001011101100",
"00010001010100111110100",
"00010001001000100000000",
"00010000111100000010011",
"00010000101111100101110",
"00010000100011001010000",
"00010000010110101110111",
"00010000001010010100110",
"00001111111101111011100",
"00001111110001100011000",
"00001111100101001011011",
"00001111011000110100110",
"00001111001100011110110",
"00001111000000001001101",
"00001110110011110101100",
"00001110100111100010000",
"00001110011011001111100",
"00001110001110111101111",
"00001110000010101101000",
"00001101110110011100110",
"00001101101010001101101",
"00001101011101111111010",
"00001101010001110001101",
"00001101000101100100111",
"00001100111001011001010",
"00001100101101001110001",
"00001100100001000011111",
"00001100010100111010011",
"00001100001000110001111",
"00001011111100101010001",
"00001011110000100011001",
"00001011100100011101001",
"00001011011000010111110",
"00001011001100010011001",
"00001011000000001111100",
"00001010110100001100101",
"00001010101000001010110",
"00001010011100001001011",
"00001010010000001001001",
"00001010000100001001011",
"00001001111000001010110",
"00001001101100001100101",
"00001001100000001111011",
"00001001010100010011001",
"00001001001000010111100",
"00001000111100011100111",
"00001000110000100010110",
"00001000100100101001101",
"00001000011000110001011",
"00001000001100111001110",
"00001000000001000011000",
"00000111110101001101001",
"00000111101001011000000",
"00000111011101100011101",
"00000111010001110000000",
"00000111000101111101010",
"00000110111010001011010",
"00000110101110011010000",
"00000110100010101001101",
"00000110010110111010001",
"00000110001011001011001",
"00000101111111011101001",
"00000101110011110000000",
"00000101101000000011011",
"00000101011100010111111",
"00000101010000101100111",
"00000101000101000010101",
"00000100111001011001010",
"00000100101101110000110",
"00000100100010001001001",
"00000100010110100010000",
"00000100001010111011110",
"00000011111111010110011",
"00000011110011110001110",
"00000011101000001101110",
"00000011011100101010100",
"00000011010001001000010",
"00000011000101100110101",
"00000010111010000101110",
"00000010101110100101110",
"00000010100011000110100",
"00000010010111100111111",
"00000010001100001010001",
"00000010000000101101001",
"00000001110101010000110",
"00000001101001110101100",
"00000001011110011010110",
"00000001010011000000101",
"00000001000111100111100",
"00000000111100001111001",
"00000000110000110111011",
"00000000100101100000011",
"00000000011010001010001",
"00000000001110110100110",
"00000000000011100000001",
"11111111110000011000010",
"11111111011001110010000",
"11111111000011001101001",
"11111110101100101001110",
"11111110010110000111111",
"11111101111111100111010",
"11111101101001001000101",
"11111101010010101011000",
"11111100111100001111001",
"11111100100101110100101",
"11111100001111011011111",
"11111011111001000100001",
"11111011100010101110000",
"11111011001100011001100",
"11111010110110000110100",
"11111010011111110101000",
"11111010001001100100110",
"11111001110011010110010",
"11111001011101001000110",
"11111001000110111101001",
"11111000110000110011000",
"11111000011010101010000",
"11111000000100100010101",
"11110111101110011100110",
"11110111011000011000001",
"11110111000010010101011",
"11110110101100010011110",
"11110110010110010011110",
"11110110000000010100111",
"11110101101010010111110",
"11110101010100011100000",
"11110100111110100001110",
"11110100101000101000101",
"11110100010010110001000",
"11110011111100111010111",
"11110011100111000110011",
"11110011010001010011011",
"11110010111011100001100",
"11110010100101110001010",
"11110010010000000010001",
"11110001111010010100110",
"11110001100100101000101",
"11110001001110111110001",
"11110000111001010100101",
"11110000100011101100110",
"11110000001110000110011",
"11101111111000100001100",
"11101111100010111101110",
"11101111001101011011101",
"11101110110111111010111",
"11101110100010011011011",
"11101110001100111101011",
"11101101110111100000111",
"11101101100010000101100",
"11101101001100101011101",
"11101100110111010011010",
"11101100100001111100001",
"11101100001100100110011",
"11101011110111010010010",
"11101011100001111111101",
"11101011001100101110000",
"11101010110111011101101",
"11101010100010001111001",
"11101010001101000001110",
"11101001110111110101111",
"11101001100010101011001",
"11101001001101100001111",
"11101000111000011010010",
"11101000100011010011101",
"11101000001110001110100",
"11100111111001001010100",
"11100111100100001000001",
"11100111001111000111001",
"11100110111010000111101",
"11100110100101001001010",
"11100110010000001100000",
"11100101111011010000101",
"11100101100110010110011",
"11100101010001011101010",
"11100100111100100101101",
"11100100100111101111100",
"11100100010010111010100",
"11100011111110000111000",
"11100011101001010101000",
"11100011010100100100000",
"11100010111111110100101",
"11100010101011000110010",
"11100010010110011001100",
"11100010000001101101110",
"11100001101101000011100",
"11100001011000011010110",
"11100001000011110011001",
"11100000101111001101000",
"11100000011010100111111",
"11100000000110000100011",
"11011111110001100010010",
"11011111011101000001010",
"11011111001000100001110",
"11011110110100000011011",
"11011110011111100110100",
"11011110001011001010101",
"11011101110110110000010",
"11011101100010010111001",
"11011101001101111111010",
"11011100111001101001000",
"11011100100101010011110",
"11011100010001000000000",
"11011011111100101101011",
"11011011101000011011111",
"11011011010100001100010",
"11011010111111111101010",
"11011010101011110000001",
"11011010010111100011110",
"11011010000011011001001",
"11011001101111001111011",
"11011001011011000111010",
"11011001000111000000011",
"11011000110010111010100",
"11011000011110110110001",
"11011000001010110010111",
"11010111110110110001001",
"11010111100010110000110",
"11010111001110110001011",
"11010110111010110011010",
"11010110100110110110100",
"11010110010010111010111",
"11010101111111000000101",
"11010101101011000111111",
"11010101010111001111111",
"11010101000011011001101",
"11010100101111100100100",
"11010100011011110000100",
"11010100000111111101111",
"11010011110100001100011",
"11010011100000011100011",
"11010011001100101101011",
"11010010111000111111100",
"11010010100101010011000",
"11010010010001101000000",
"11010001111101111110000",
"11010001101010010101100",
"11010001010110101101110",
"11010001000011000111110",
"11010000101111100010110",
"11010000011011111111000",
"11010000001000011100100",
"11001111110100111011010",
"11001111100001011011000",
"11001111001101111100100",
"11001110111010011110110",
"11001110100111000010011",
"11001110010011100111001",
"11001110000000001101010",
"11001101101100110100100",
"11001101011001011101010",
"11001101000110000111000",
"11001100110010110001110",
"11001100011111011110000",
"11001100001100001011010",
"11001011111000111010000",
"11001011100101101001110",
"11001011010010011011000",
"11001010111111001101010",
"11001010101100000000100",
"11001010011000110101010",
"11001010000101101011001",
"11001001110010100010000",
"11001001011111011010010",
"11001001001100010011101",
"11001000111001001110011",
"11001000100110001010001",
"11001000010011000111000",
"11001000000000000101011",
"11000111101101000100101",
"11000111011010000101011",
"11000111000111000111010",
"11000110110100001010001",
"11000110100001001110011",
"11000110001110010011101",
"11000101111011011010000",
"11000101101000100001110",
"11000101010101101010101",
"11000101000010110100111",
"11000100101111111111110",
"11000100011101001100100",
"11000100001010011001111",
"11000011110111101000101",
"11000011100100111000100",
"11000011010010001001101",
"11000010111111011011111",
"11000010101100101111010",
"11000010011010000011101",
"11000010000111011001011",
"11000001110100110000100",
"11000001100010001000011",
"11000001001111100001100",
"11000000111100111011111",
"11000000101010010111100",
"11000000010111110100001",
"11000000000101010001111",
"10111111110010110000110",
"10111111100000010000111",
"10111111001101110010000",
"10111110111011010100101",
"10111110101000110111111",
"10111110010110011100111",
"10111110000100000010101",
"10111101110001101001101",
"10111101011111010001100",
"10111101001100111010111",
"10111100111010100101001",
"10111100101000010000101",
"10111100010101111101010",
"10111100000011101011010",
"10111011110001011001111",
"10111011011111001001111",
"10111011001100111010111",
"10111010111010101101011",
"10111010101000100000110",
"10111010010110010101010",
"10111010000100001010110",
"10111001110010000001101",
"10111001011111111001100",
"10111001001101110010011",
"10111000111011101100011",
"10111000101001100111110",
"10111000010111100100000",
"10111000000101100001011",
"10110111110011011111110",
"10110111100001011111100",
"10110111001111100000010",
"10110110111101100010000",
"10110110101011100101001",
"10110110011001101001000",
"10110110000111101110001",
"10110101110101110100011",
"10110101100011111011111",
"10110101010010000100001",
"10110101000000001101110",
"10110100101110011000010",
"10110100011100100100010",
"10110100001010110000111",
"10110011111000111110111",
"10110011100111001101110",
"10110011010101011101110",
"10110011000011101111001",
"10110010110010000001001",
"10110010100000010100100",
"10110010001110101000111",
"10110001111100111110010",
"10110001101011010101000",
"10110001011001101100110",
"10110001001000000101100",
"10110000110110011111010",
"10110000100100111010000",
"10110000010011010101110",
"10110000000001110010111",
"10101111110000010000111",
"10101111011110110000000",
"10101111001101010000001",
"10101110111011110001100",
"10101110101010010011101",
"10101110011000110111001",
"10101110000111011011100",
"10101101110110000001000",
"10101101100100100111110",
"10101101010011001111010",
"10101101000001111000000",
"10101100110000100001110",
"10101100011111001100100",
"10101100001101111000010",
"10101011111100100101000",
"10101011101011010011001",
"10101011011010000001111",
"10101011001000110001111",
"10101010110111100011000",
"10101010100110010101000",
"10101010010101001000011",
"10101010000011111100011",
"10101001110010110001110",
"10101001100001100111110",
"10101001010000011111001",
"10101000111111010111011",
"10101000101110010000110",
"10101000011101001011011",
"10101000001100000110101",
"10100111111011000011010",
"10100111101010000000100",
"10100111011000111111000",
"10100111000111111110101",
"10100110110110111111001",
"10100110100110000000101",
"10100110010101000011100",
"10100110000100000110111",
"10100101110011001011110",
"10100101100010010001001",
"10100101010001010111111",
"10100101000000011111101",
"10100100101111101000011",
"10100100011110110010000",
"10100100001101111100101",
"10100011111101001000011",
"10100011101100010101010",
"10100011011011100010111",
"10100011001010110001110",
"10100010111010000001101",
"10100010101001010010001",
"10100010011000100011111",
"10100010000111110110110",
"10100001110111001010100",
"10100001100110011111100",
"10100001010101110101010",
"10100001000101001011111",
"10100000110100100011100",
"10100000100011111100100",
"10100000010011010110000",
"10100000000010110000111",
"10011111110010001100110",
"10011111100001101001100",
"10011111010001000111000",
"10011111000000100101110",
"10011110110000000101011",
"10011110011111100110000",
"10011110001111000111101",
"10011101111110101010010",
"10011101101110001110001",
"10011101011101110010101",
"10011101001101011000001",
"10011100111100111110111",
"10011100101100100110010",
"10011100011100001110101",
"10011100001011111000010",
"10011011111011100010100",
"10011011101011001110001",
"10011011011010111010101",
"10011011001010100111110",
"10011010111010010110001",
"10011010101010000101100",
"10011010011001110101100",
"10011010001001100110111",
"10011001111001011001000",
"10011001101001001100010",
"10011001011001000000011",
"10011001001000110101100",
"10011000111000101011100",
"10011000101000100010010",
"10011000011000011010001",
"10011000001000010011000",
"10010111111000001100111",
"10010111101000000111110",
"10010111011000000011100",
"10010111001000000000001",
"10010110110111111101110",
"10010110100111111100011",
"10010110010111111011111",
"10010110000111111100011",
"10010101110111111101110",
"10010101101000000000001",
"10010101011000000011011",
"10010101001000000111101",
"10010100111000001100111",
"10010100101000010011000",
"10010100011000011010001",
"10010100001000100010001",
"10010011111000101011000",
"10010011101000110100111",
"10010011011000111111110",
"10010011001001001011100",
"10010010111001011000010",
"10010010101001100101100",
"10010010011001110100001",
"10010010001010000011101",
"10010001111010010100001",
"10010001101010100101001",
"10010001011010110111100",
"10010001001011001010110",
"10010000111011011110101",
"10010000101011110011110",
"10010000011100001001011",
"10010000001100100000011",
"10001111111100111000000",
"10001111101101010000111",
"10001111011101101010010",
"10001111001110000100101",
"10001110111110100000000",
"10001110101110111100010",
"10001110011111011001110",
"10001110001111110111111",
"10001110000000010110111",
"10001101110000110110110",
"10001101100001010111011",
"10001101010001111001001",
"10001101000010011011111",
"10001100110010111111100",
"10001100100011100011110",
"10001100010100001001010",
"10001100000100101111011",
"10001011110101010110101",
"10001011100101111110101",
"10001011010110100111100",
"10001011000111010001010",
"10001010110111111100000",
"10001010101000100111101",
"10001010011001010100001",
"10001010001010000001100",
"10001001111010101111111",
"10001001101011011110111",
"10001001011100001111001",
"10001001001100111111111",
"10001000111101110001101",
"10001000101110100100101",
"10001000011111011000001",
"10001000010000001100101",
"10001000000001000010000",
"10000111110001111000010",
"10000111100010101111001",
"10000111010011100111010",
"10000111000100100000000",
"10000110110101011001111",
"10000110100110010100011",
"10000110010111001111111",
"10000110001000001100001",
"10000101111001001001011",
"10000101101010000111101",
"10000101011011000110101",
"10000101001100000110011",
"10000100111101000111010",
"10000100101110001000101",
"10000100011111001011000",
"10000100010000001110011",
"10000100000001010010100",
"10000011110010010111101",
"10000011100011011101010",
"10000011010100100100001",
"10000011000101101011101",
"10000010110110110100000",
"10000010100111111101101",
"10000010011001000111100",
"10000010001010010010101",
"10000001111011011110101",
"10000001101100101011001",
"10000001011101111000111",
"10000001001111000111010",
"10000001000000010110100",
"10000000110001100110110",
"10000000100010110111110",
"10000000010100001001011",
"10000000000101011100000",
"01111111110110101111110",
"01111111101000000100000",
"01111111011001011001010",
"01111111001010101111000",
"01111110111100000110000",
"01111110101101011101101",
"01111110011110110110011",
"01111110010000001111110",
"01111110000001101010000",
"01111101110011000100111",
"01111101100100100000111",
"01111101010101111101100",
"01111101000111011011000",
"01111100111000111001100",
"01111100101010011000110",
"01111100011011111000111",
"01111100001101011001101",
"01111011111110111011010",
"01111011110000011101110",
"01111011100010000001010",
"01111011010011100101100",
"01111011000101001010011",
"01111010110110110000011",
"01111010101000010111000",
"01111010011001111110100",
"01111010001011100110101",
"01111001111101001111111",
"01111001101110111001110",
"01111001100000100100100",
"01111001010010010000001",
"01111001000011111100010",
"01111000110101101001101",
"01111000100111010111100",
"01111000011001000110011",
"01111000001010110110000",
"01110111111100100110011",
"01110111101110010111100",
"01110111100000001001110",
"01110111010001111100011",
"01110111000011110000001",
"01110110110101100100110",
"01110110100111011010000",
"01110110011001010000000",
"01110110001011000110101",
"01110101111100111110100",
"01110101101110110110111",
"01110101100000110000001",
"01110101010010101010010",
"01110101000100100101010",
"01110100110110100000111",
"01110100101000011101010",
"01110100011010011010101",
"01110100001100011000100",
"01110011111110010111100",
"01110011110000010111001",
"01110011100010010111101",
"01110011010100011000101",
"01110011000110011010100",
"01110010111000011101010",
"01110010101010100000111",
"01110010011100100101011",
"01110010001110101010100",
"01110010000000110000011",
"01110001110010110111001",
"01110001100100111110100",
"01110001010111000111000",
"01110001001001010000001",
"01110000111011011001110",
"01110000101101100100100",
"01110000011111101111111",
"01110000010001111100000",
"01110000000100001001001",
"01101111110110010110110",
"01101111101000100101001",
"01101111011010110100100",
"01101111001101000100011",
"01101110111111010101001",
"01101110110001100110110",
"01101110100011111001010",
"01101110010110001100010",
"01101110001000100000001",
"01101101111010110100110",
"01101101101101001010011",
"01101101011111100000100",
"01101101010001110111100",
"01101101000100001111010",
"01101100110110100111110",
"01101100101001000000111",
"01101100011011011011000",
"01101100001101110101101",
"01101100000000010001001",
"01101011110010101101100",
"01101011100101001010011",
"01101011010111101000011",
"01101011001010000111000",
"01101010111100100110001",
"01101010101111000110001",
"01101010100001100110111",
"01101010010100001000101",
"01101010000110101010110",
"01101001111001001101111",
"01101001101011110001110",
"01101001011110010110010",
"01101001010000111011100",
"01101001000011100001101",
"01101000110110001000101",
"01101000101000110000001",
"01101000011011011000010",
"01101000001110000001011",
"01101000000000101011001",
"01100111110011010101110",
"01100111100110000000111",
"01100111011000101100111",
"01100111001011011001110",
"01100110111110000111000",
"01100110110000110101010",
"01100110100011100100010",
"01100110010110010011111",
"01100110001001000100010",
"01100101111011110101100",
"01100101101110100111101",
"01100101100001011001111",
"01100101010100001101011",
"01100101000111000001011",
"01100100111001110110001",
"01100100101100101011111",
"01100100011111100010000",
"01100100010010011001001",
"01100100000101010000111",
"01100011111000001001011",
"01100011101011000010100",
"01100011011101111100011",
"01100011010000110110111",
"01100011000011110010011",
"01100010110110101110010",
"01100010101001101011001",
"01100010011100101000110",
"01100010001111100110111",
"01100010000010100101111",
"01100001110101100101011",
"01100001101000100101110",
"01100001011011100110111",
"01100001001110101000111",
"01100001000001101011011",
"01100000110100101110100",
"01100000100111110010011",
"01100000011010110111000",
"01100000001101111100100",
"01100000000001000010101",
"01011111110100001001010",
"01011111100111010000111",
"01011111011010011001001",
"01011111001101100001111",
"01011111000000101011100",
"01011110110011110101111",
"01011110100111000000110",
"01011110011010001100100",
"01011110001101011001001",
"01011110000000100110010",
"01011101110011110011111",
"01011101100111000010100",
"01011101011010010001110",
"01011101001101100001101",
"01011101000000110010001",
"01011100110100000011101",
"01011100100111010101100",
"01011100011010101000010",
"01011100001101111011111",
"01011100000001001111111",
"01011011110100100100100",
"01011011100111111010010",
"01011011011011010000010",
"01011011001110100111010",
"01011011000001111110111",
"01011010110101010110111",
"01011010101000101111110",
"01011010011100001001100",
"01011010001111100011110",
"01011010000010111110110",
"01011001110110011010101",
"01011001101001110111000",
"01011001011101010011111",
"01011001010000110001101",
"01011001000100010000001",
"01011000110111101111001",
"01011000101011001111000",
"01011000011110101111011",
"01011000010010010000100",
"01011000000101110010100",
"01010111111001010100111",
"01010111101100110111111",
"01010111100000011100000",
"01010111010100000000011",
"01010111000111100101110",
"01010110111011001011011",
"01010110101110110010001",
"01010110100010011001010",
"01010110010110000001000",
"01010110001001101001101",
"01010101111101010011000",
"01010101110000111100111",
"01010101100100100111100",
"01010101011000010010101",
"01010101001011111110101",
"01010100111111101011001",
"01010100110011011000011",
"01010100100111000110010",
"01010100011010110100110",
"01010100001110100011111",
"01010100000010010011110",
"01010011110110000100100",
"01010011101001110101110",
"01010011011101100111011",
"01010011010001011001111",
"01010011000101001101010",
"01010010111001000001000",
"01010010101100110101101",
"01010010100000101010110",
"01010010010100100000011",
"01010010001000010111000",
"01010001111100001110000",
"01010001110000000110000",
"01010001100011111110001",
"01010001010111110111100",
"01010001001011110001000",
"01010000111111101011100",
"01010000110011100110011",
"01010000100111100010010",
"01010000011011011110101",
"01010000001111011011100",
"01010000000011011001001",
"01001111110111010111011",
"01001111101011010110010",
"01001111011111010101110",
"01001111010011010110000",
"01001111000111010110110",
"01001110111011011000010",
"01001110101111011010101",
"01001110100011011101001",
"01001110010111100000110",
"01001110001011100100101",
"01001101111111101001100",
"01001101110011101110111",
"01001101100111110100110",
"01001101011011111011011",
"01001101010000000010101",
"01001101000100001010100",
"01001100111000010011000",
"01001100101100011100000",
"01001100100000100110000",
"01001100010100110000001",
"01001100001000111011001",
"01001011111101000111000",
"01001011110001010011010",
"01001011100101100000010",
"01001011011001101101111",
"01001011001101111011111",
"01001011000010001010110",
"01001010110110011010010",
"01001010101010101010011",
"01001010011110111011000",
"01001010010011001100011",
"01001010000111011110001",
"01001001111011110000110",
"01001001110000000011111",
"01001001100100010111111",
"01001001011000101100010",
"01001001001101000001011",
"01001001000001010111000",
"01001000110101101101011",
"01001000101010000100011",
"01001000011110011011110",
"01001000010010110011111",
"01001000000111001100101",
"01000111111011100110000",
"01000111110000000000000",
"01000111100100011010101",
"01000111011000110101110",
"01000111001101010001110",
"01000111000001101110010",
"01000110110110001011011",
"01000110101010101001001",
"01000110011111000111010",
"01000110010011100110010",
"01000110001000000101101",
"01000101111100100101111",
"01000101110001000110100",
"01000101100101100111110",
"01000101011010001001101",
"01000101001110101100011",
"01000101000011001111100",
"01000100110111110011001",
"01000100101100010111101",
"01000100100000111100100",
"01000100010101100010010",
"01000100001010001000011",
"01000011111110101111000",
"01000011110011010110011",
"01000011100111111110010",
"01000011011100100110111",
"01000011010001010000001",
"01000011000101111010000",
"01000010111010100100011",
"01000010101111001111001",
"01000010100011111010110",
"01000010011000100110111",
"01000010001101010011110",
"01000010000010000001000",
"01000001110110101110111",
"01000001101011011101011",
"01000001100000001100100",
"01000001010100111100010",
"01000001001001101100100",
"01000000111110011101100",
"01000000110011001110110",
"01000000101000000001000",
"01000000011100110011100",
"01000000010001100111000",
"01000000000110011010101",
"00111111111011001111001",
"00111111110000000100000",
"00111111100100111001110",
"00111111011001101111111",
"00111111001110100110100",
"00111111000011011101111",
"00111110111000010110000",
"00111110101101001110010",
"00111110100010000111011",
"00111110010111000001001",
"00111110001011111011100",
"00111110000000110110010",
"00111101110101110001100",
"00111101101010101101100",
"00111101011111101010010",
"00111101010100100111001",
"00111101001001100100110",
"00111100111110100011010",
"00111100110011100010001",
"00111100101000100001100",
"00111100011101100001101",
"00111100010010100010010",
"00111100000111100011010",
"00111011111100100101000",
"00111011110001100111010",
"00111011100110101010000",
"00111011011011101101100",
"00111011010000110001100",
"00111011000101110110001",
"00111010111010111011010",
"00111010110000000000111",
"00111010100101000111010",
"00111010011010001110001",
"00111010001111010101011",
"00111010000100011101100",
"00111001111001100110000",
"00111001101110101111010",
"00111001100011111000111",
"00111001011001000011001",
"00111001001110001101110",
"00111001000011011001001",
"00111000111000100101010",
"00111000101101110001100",
"00111000100010111110101",
"00111000011000001100001",
"00111000001101011010011",
"00111000000010101001000",
"00110111110111111000010",
"00110111101101001000001",
"00110111100010011000100",
"00110111010111101001011",
"00110111001100111010111",
"00110111000010001100111",
"00110110110111011111101",
"00110110101100110010101",
"00110110100010000110010",
"00110110010111011010110",
"00110110001100101111101",
"00110110000010000100111",
"00110101110111011010110",
"00110101101100110001010",
"00110101100010001000010",
"00110101010111011111101",
"00110101001100110111111",
"00110101000010010000100",
"00110100110111101001101",
"00110100101101000011011",
"00110100100010011101101",
"00110100010111111000101",
"00110100001101010011111",
"00110100000010101111110",
"00110011111000001100011",
"00110011101101101001010",
"00110011100011000110110",
"00110011011000100100110",
"00110011001110000011100",
"00110011000011100010110",
"00110010111001000010011",
"00110010101110100010110",
"00110010100100000011010",
"00110010011001100100111",
"00110010001111000110101",
"00110010000100101001000",
"00110001111010001100000",
"00110001101111101111010",
"00110001100101010011011",
"00110001011010110111111",
"00110001010000011100111",
"00110001000110000010101",
"00110000111011101000110",
"00110000110001001111011",
"00110000100110110110100",
"00110000011100011110010",
"00110000010010000110100",
"00110000000111101111011",
"00101111111101011000100",
"00101111110011000010011",
"00101111101000101101000",
"00101111011110010111110",
"00101111010100000011010",
"00101111001001101111001",
"00101110111111011011110",
"00101110110101001000101",
"00101110101010110110001",
"00101110100000100100011",
"00101110010110010010110",
"00101110001100000001111",
"00101110000001110001100",
"00101101110111100001110",
"00101101101101010010010",
"00101101100011000011100",
"00101101011000110101001",
"00101101001110100111100",
"00101101000100011010010",
"00101100111010001101100",
"00101100110000000001001",
"00101100100101110101101",
"00101100011011101010011",
"00101100010001011111110",
"00101100000111010101100",
"00101011111101001011111",
"00101011110011000010110",
"00101011101000111010001",
"00101011011110110010001",
"00101011010100101010101",
"00101011001010100011100",
"00101011000000011100111",
"00101010110110010111000",
"00101010101100010001010",
"00101010100010001100100",
"00101010011000000111111",
"00101010001110000100000",
"00101010000100000000010",
"00101001111001111101100",
"00101001101111111010111",
"00101001100101111001000",
"00101001011011110111011",
"00101001010001110110101",
"00101001000111110110000",
"00101000111101110110010",
"00101000110011110110110",
"00101000101001110111110",
"00101000011111111001010",
"00101000010101111011100",
"00101000001011111110000",
"00101000000010000001001",
"00100111111000000100101",
"00100111101110001000110",
"00100111100100001101011",
"00100111011010010010011",
"00100111010000010111111",
"00100111000110011110001",
"00100110111100100100100",
"00100110110010101011100",
"00100110101000110011010",
"00100110011110111011010",
"00100110010101000011111",
"00100110001011001100111",
"00100110000001010110011",
"00100101110111100000101",
"00100101101101101011000",
"00100101100011110110000",
"00100101011010000001100",
"00100101010000001101110",
"00100101000110011010000",
"00100100111100100111001",
"00100100110010110100101",
"00100100101001000010100",
"00100100011111010001001",
"00100100010101100000001",
"00100100001011101111011",
"00100100000001111111100",
"00100011111000001111111",
"00100011101110100000111",
"00100011100100110010001",
"00100011011011000100000",
"00100011010001010110101",
"00100011000111101001011",
"00100010111101111100110",
"00100010110100010000101",
"00100010101010100101000",
"00100010100000111001101",
"00100010010111001110111",
"00100010001101100100101",
"00100010000011111011000",
"00100001111010010001101",
"00100001110000101000110",
"00100001100111000000101",
"00100001011101011000111",
"00100001010011110001100",
"00100001001010001010101",
"00100001000000100100001",
"00100000110110111110011",
"00100000101101011000110",
"00100000100011110011110",
"00100000011010001111010",
"00100000010000101011011",
"00100000000111000111110",
"00011111111101100100110",
"00011111110100000010010",
"00011111101010100000001",
"00011111100000111110011",
"00011111010111011101011",
"00011111001101111100100",
"00011111000100011100011",
"00011110111010111100100",
"00011110110001011101010",
"00011110100111111110101",
"00011110011110100000001",
"00011110010101000010010",
"00011110001011100100111",
"00011110000010000111111",
"00011101111000101011101",
"00011101101111001111100",
"00011101100101110100001",
"00011101011100011001000",
"00011101010010111110100",
"00011101001001100100010",
"00011101000000001010100",
"00011100110110110001011",
"00011100101101011000110",
"00011100100100000000100",
"00011100011010101000110",
"00011100010001010001010",
"00011100000111111010010",
"00011011111110100100000",
"00011011110101001110001",
"00011011101011111000101",
"00011011100010100011101",
"00011011011001001110111",
"00011011001111111010110",
"00011011000110100111001",
"00011010111101010100000",
"00011010110100000001010",
"00011010101010101111000",
"00011010100001011101001",
"00011010011000001011101",
"00011010001110111010111",
"00011010000101101010100",
"00011001111100011010010",
"00011001110011001011000",
"00011001101001111011111",
"00011001100000101101001",
"00011001010111011111000",
"00011001001110010001001",
"00011001000101000011111",
"00011000111011110111001",
"00011000110010101010110",
"00011000101001011110110",
"00011000100000010011011",
"00011000010111001000010",
"00011000001101111101110",
"00011000000100110011110",
"00010111111011101010000",
"00010111110010100000110",
"00010111101001010111111",
"00010111100000001111100",
"00010111010111000111110",
"00010111001110000000011",
"00010111000100111001001",
"00010110111011110010101",
"00010110110010101100100",
"00010110101001100111001",
"00010110100000100001110",
"00010110010111011101001",
"00010110001110011000101",
"00010110000101010100111",
"00010101111100010001011",
"00010101110011001110011",
"00010101101010001011110",
"00010101100001001001101",
"00010101011000001000001",
"00010101001111000110110",
"00010101000110000110000",
"00010100111101000101110",
"00010100110100000101111",
"00010100101011000110011",
"00010100100010000111010",
"00010100011001001000101",
"00010100010000001010100",
"00010100000111001100110",
"00010011111110001111100",
"00010011110101010010110",
"00010011101100010110010",
"00010011100011011010011",
"00010011011010011110110",
"00010011010001100011100",
"00010011001000101000110",
"00010010111111101110101",
"00010010110110110100110",
"00010010101101111011011",
"00010010100101000010100",
"00010010011100001010000",
"00010010010011010001111",
"00010010001010011010010",
"00010010000001100010111",
"00010001111000101100010",
"00010001101111110101110",
"00010001100111000000000",
"00010001011110001010010",
"00010001010101010101010",
"00010001001100100000101",
"00010001000011101100011",
"00010000111010111000100",
"00010000110010000101001",
"00010000101001010010011",
"00010000100000011111110",
"00010000010111101101100",
"00010000001110111100000",
"00010000000110001010110",
"00001111111101011001110",
"00001111110100101001011",
"00001111101011111001011",
"00001111100011001001111",
"00001111011010011010111",
"00001111010001101100001",
"00001111001000111101110",
"00001111000000010000000",
"00001110110111100010011",
"00001110101110110101100",
"00001110100110001000110",
"00001110011101011100100",
"00001110010100110000111",
"00001110001100000101100",
"00001110000011011010100",
"00001101111010110000000",
"00001101110010000101110",
"00001101101001011100010",
"00001101100000110010111",
"00001101011000001010000",
"00001101001111100001101",
"00001101000110111001100",
"00001100111110010001111",
"00001100110101101010110",
"00001100101101000100000",
"00001100100100011101110",
"00001100011011110111110",
"00001100010011010010001",
"00001100001010101101000",
"00001100000010001000010",
"00001011111001100011111",
"00001011110001000000001",
"00001011101000011100100",
"00001011011111111001010",
"00001011010111010110110",
"00001011001110110100101",
"00001011000110010010100",
"00001010111101110001001",
"00001010110101010000001",
"00001010101100101111100",
"00001010100100001111011",
"00001010011011101111100",
"00001010010011010000001",
"00001010001010110001000",
"00001010000010010010011",
"00001001111001110100001",
"00001001110001010110100",
"00001001101000111001000",
"00001001100000011100000",
"00001001010111111111100",
"00001001001111100011010",
"00001001000111000111100",
"00001000111110101100010",
"00001000110110010001001",
"00001000101101110110101",
"00001000100101011100100",
"00001000011101000010110",
"00001000010100101001011",
"00001000001100010000100",
"00001000000011110111111",
"00000111111011011111110",
"00000111110011000111111",
"00000111101010110000100",
"00000111100010011001100",
"00000111011010000010111",
"00000111010001101100101",
"00000111001001010111000",
"00000111000001000001100",
"00000110111000101100011",
"00000110110000011000000",
"00000110101000000011101",
"00000110011111110000000",
"00000110010111011100011",
"00000110001111001001100",
"00000110000110110110111",
"00000101111110100100100",
"00000101110110010010110",
"00000101101110000001011",
"00000101100101110000011",
"00000101011101011111100",
"00000101010101001111010",
"00000101001100111111100",
"00000101000100110000000",
"00000100111100100000111",
"00000100110100010010010",
"00000100101100000011111",
"00000100100011110110000",
"00000100011011101000011",
"00000100010011011011010",
"00000100001011001110011",
"00000100000011000010000",
"00000011111010110110000",
"00000011110010101010011",
"00000011101010011111011",
"00000011100010010100011",
"00000011011010001001111",
"00000011010001111111110",
"00000011001001110110000",
"00000011000001101100111",
"00000010111001100011111",
"00000010110001011011011",
"00000010101001010011011",
"00000010100001001011100",
"00000010011001000100000",
"00000010010000111101001",
"00000010001000110110100",
"00000010000000110000011",
"00000001111000101010011",
"00000001110000100100111",
"00000001101000011111111",
"00000001100000011011000",
"00000001011000010110111",
"00000001010000010010110",
"00000001001000001111011",
"00000001000000001100000",
"00000000111000001001011",
"00000000110000000110110",
"00000000101000000100111",
"00000000100000000011000",
"00000000011000000001111",
"00000000010000000000110",
"00000000001000000000011");

begin

  data<=rom1(conv_integer(addr));
  data2<=rom2(conv_integer(addr));

  end VHDL;
