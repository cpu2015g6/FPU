library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.STD_LOGIC_ARITH.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity fputop is
  port(MCLK1: in std_logic;
       RS_TX: out std_logic);
  end fputop;

architecture VHDL of fputop is

component fadd
  port(clk: in std_logic;
       op1, op2:  in std_logic_vector(31 downto 0);
       ans:       out std_logic_vector(31 downto 0) := x"00000000"
       );
end component;

component u232c
  generic (wtime: std_logic_vector(15 downto 0) := x"1ADB");
  Port ( clk  : in  STD_LOGIC;
         data : in  STD_LOGIC_VECTOR (7 downto 0);
         go   : in  STD_LOGIC;
         busy : out STD_LOGIC;
         tx   : out STD_LOGIC);
end component;

  signal clk,iclk: std_logic;
  type rom_t is array(0 to 497) of std_logic_vector(31 downto 0);
  constant rom: rom_t := ("00111111100000000000000000000000",
"00111111100000000000000000000000",
"01000000000000000000000000000000",
"10111111100000000000000000000000",
"10111111100000000000000000000000",
"11000000000000000000000000000000",
"00001011111111111111111111111111",
"10001100000000000000000000000000",
"10000000010000000000000000000000",
"00001011111111111111111111111110",
"10001100000000000000000000000000",
"10000000100000000000000000000000",
"00001100011111111111111111111111",
"10001100100000000000000000000000",
"10000000100000000000000000000000",
"11111101010010010100110010111110",
"01111001000111011100100001010111",
"11111101010010001010111011110110",
"01111001000111011100100001010111",
"11111101010010010100110010111110",
"11111101010010001010111011110110",
"00000011101111000000110100101101",
"10010001001001111001110101011000",
"10010001001001111001110101011000",
"10010001001001111001110101011000",
"00000011101111000000110100101101",
"10010001001001111001110101011000",
"00011000110000111011011100111110",
"10010011011101010000010001101110",
"00011000110000111001100010011101",
"10010011011101010000010001101110",
"00011000110000111011011100111110",
"00011000110000111001100010011101",
"11010100101011100100000011100100",
"11011000110100010110011100001000",
"11011000110100100001010101001001",
"11011000110100010110011100001000",
"11010100101011100100000011100100",
"11011000110100100001010101001001",
"01110101010010110000010001010100",
"10000100010001001100001101111001",
"01110101010010110000010001010100",
"10000100010001001100001101111001",
"01110101010010110000010001010100",
"01110101010010110000010001010100",
"10101101011111100011010010110111",
"00111000000100001010100010011101",
"00111000000100001010100010011001",
"00111000000100001010100010011101",
"10101101011111100011010010110111",
"00111000000100001010100010011001",
"00011000011010000101000001010000",
"00011100011000101010001000011001",
"00011100011000111000101001101001",
"00011100011000101010001000011001",
"00011000011010000101000001010000",
"00011100011000111000101001101001",
"10000011111010100000011110001001",
"10001001110110100010110101110100",
"10001001110110100011110000010100",
"10001001110110100010110101110100",
"10000011111010100000011110001001",
"10001001110110100011110000010100",
"00001101010000111111111000010101",
"10000010010001100110011001111011",
"00001101010000111111111000010010",
"10000010010001100110011001111011",
"00001101010000111111111000010101",
"00001101010000111111111000010010",
"11000100011011101001011011100111",
"11001110110011110110101100101001",
"11001110110011110110101100110000",
"11001110110011110110101100101001",
"11000100011011101001011011100111",
"11001110110011110110101100110000",
"00010011000010100101100110000100",
"10001000011000110010110010101100",
"00010011000010100101100110000000",
"10001000011000110010110010101100",
"00010011000010100101100110000100",
"00010011000010100101100110000000",
"10001000010110000001100000100110",
"11111101110111111011011011010000",
"11111101110111111011011011010000",
"11111101110111111011011011010000",
"10001000010110000001100000100110",
"11111101110111111011011011010000",
"10111001100111110000000001110000",
"10101010110011101010011001001101",
"10111001100111110000000001110000",
"10101010110011101010011001001101",
"10111001100111110000000001110000",
"10111001100111110000000001110000",
"10101001001101000000100110010110",
"10101000011010010000000001000000",
"10101001011011100100100110100110",
"10101000011010010000000001000000",
"10101001001101000000100110010110",
"10101001011011100100100110100110",
"00110110011001000111101000101001",
"00111010000101011011110111001010",
"00111010000101101010001001000100",
"00111010000101011011110111001010",
"00110110011001000111101000101001",
"00111010000101101010001001000100",
"01111110110100000111001000000010",
"01110011111100001111101011000011",
"01111110110100000111001000000110",
"01110011111100001111101011000011",
"01111110110100000111001000000010",
"01111110110100000111001000000110",
"10010100101000010011101011010000",
"00010111100111000000101000100100",
"00010111100110011000010100111001",
"00010111100111000000101000100100",
"10010100101000010011101011010000",
"00010111100110011000010100111001",
"10110011011101011111011110110111",
"00111010000111110010110010110011",
"00111010000111110010100011011011",
"00111010000111110010110010110011",
"10110011011101011111011110110111",
"00111010000111110010100011011011",
"10010000001000110110011011010000",
"10011010111101111111001100101100",
"10011010111101111111001100110001",
"10011010111101111111001100101100",
"10010000001000110110011011010000",
"10011010111101111111001100110001",
"00100110100011111011000110011110",
"10101000100100010100011001111001",
"10101000100010000100101101011111",
"10101000100100010100011001111001",
"00100110100011111011000110011110",
"10101000100010000100101101011111",
"00010000011111010000011000011100",
"00001111101001010100011011001100",
"00010000101001111101010011000001",
"00001111101001010100011011001100",
"00010000011111010000011000011100",
"00010000101001111101010011000001",
"10010111111001000101111100110001",
"00100011010100011110011000110111",
"00100011010100011110011000110101",
"00100011010100011110011000110111",
"10010111111001000101111100110001",
"00100011010100011110011000110101",
"01100101011100101111111010110111",
"11011011110110100011100011111111",
"01100101011100101111111010011100",
"11011011110110100011100011111111",
"01100101011100101111111010110111",
"01100101011100101111111010011100",
"00100000100110001010111011010111",
"10011100011011010110101100110101",
"00100000100110000011100000100001",
"10011100011011010110101100110101",
"00100000100110001010111011010111",
"00100000100110000011100000100001",
"00110011101011110111110011010000",
"10100110101001001000001001100100",
"00110011101011110111110011010000",
"10100110101001001000001001100100",
"00110011101011110111110011010000",
"00110011101011110111110011010000",
"00110001011001000110010111110000",
"00101110011001011101011011110000",
"00110001011001111111110101001100",
"00101110011001011101011011110000",
"00110001011001000110010111110000",
"00110001011001111111110101001100",
"10101011110100111101000111100111",
"10101011000010100110101010001000",
"10101100000011001000001110010110",
"10101011000010100110101010001000",
"10101011110100111101000111100111",
"10101100000011001000001110010110",
"01100011110000101011100011011000",
"01100000001010110000000110101110",
"01100011110001000000111011011011",
"01100000001010110000000110101110",
"01100011110000101011100011011000",
"01100011110001000000111011011011",
"00101101110010010010111001010100",
"00110000001110110101011101001101",
"00110000010000011010000011000000",
"00110000001110110101011101001101",
"00101101110010010010111001010100",
"00110000010000011010000011000000",
"00010110001100011101011110101001",
"00010011011011101110000010110101",
"00010110001101011001001100101100",
"00010011011011101110000010110101",
"00010110001100011101011110101001",
"00010110001101011001001100101100",
"00111010111010110010000110110001",
"11000110111111110011010111011010",
"11000110111111110011010111011001",
"11000110111111110011010111011010",
"00111010111010110010000110110001",
"11000110111111110011010111011001",
"00100010011111100111110000000000",
"00011101111110110011011101010111",
"00100010011111101111100110011100",
"00011101111110110011011101010111",
"00100010011111100111110000000000",
"00100010011111101111100110011100",
"00110001110110001100100000110011",
"11000000100101110010110001110100",
"11000000100101110010110001110100",
"11000000100101110010110001110100",
"00110001110110001100100000110011",
"11000000100101110010110001110100",
"11101110011100110110100111010011",
"01110000100111011011110101111110",
"01110000100101100010001000101111",
"01110000100111011011110101111110",
"11101110011100110110100111010011",
"01110000100101100010001000101111",
"01001111000001000111101100000011",
"01011100110011001011111011000001",
"01011100110011001011111011000001",
"01011100110011001011111011000001",
"01001111000001000111101100000011",
"01011100110011001011111011000001",
"00001000000011010111000000111001",
"00010100001111011100111001011000",
"00010100001111011100111001011001",
"00010100001111011100111001011000",
"00001000000011010111000000111001",
"00010100001111011100111001011001",
"10000101101111010100100010110010",
"10000001110100100110110010000100",
"10000101101111100001101100011111",
"10000001110100100110110010000100",
"10000101101111010100100010110010",
"10000101101111100001101100011111",
"10010001110001111001111100101100",
"10011111110100001010110101111110",
"10011111110100001010110101111110",
"10011111110100001010110101111110",
"10010001110001111001111100101100",
"10011111110100001010110101111110",
"01011010010111010011011101110111",
"11100100110011101111110111101111",
"11100100110011101111110111101000",
"11100100110011101111110111101111",
"01011010010111010011011101110111",
"11100100110011101111110111101000",
"10011001110010111110110011110000",
"00001101100111101001011000110001",
"10011001110010111110110011101111",
"00001101100111101001011000110001",
"10011001110010111110110011110000",
"10011001110010111110110011101111",
"01010010011000001010100001010111",
"11010110100010100110001010000111",
"11010110100010011111001000110011",
"11010110100010100110001010000111",
"01010010011000001010100001010111",
"11010110100010011111001000110011",
"00011001001011111011100000001001",
"00100111110110101000100101101011",
"00100111110110101000100101101011",
"00100111110110101000100101101011",
"00011001001011111011100000001001",
"00100111110110101000100101101011",
"00011001111000010010111001101101",
"00101001011010100011001010101000",
"00101001011010100011001010101000",
"00101001011010100011001010101000",
"00011001111000010010111001101101",
"00101001011010100011001010101000",
"01110000110101100110110100010010",
"01111010010101001011011100100011",
"01111010010101001011011100111110",
"01111010010101001011011100100011",
"01110000110101100110110100010010",
"01111010010101001011011100111110",
"10100100011000110011011011011001",
"00011110100111100110000110111010",
"10100100011000110010001100001101",
"00011110100111100110000110111010",
"10100100011000110011011011011001",
"10100100011000110010001100001101",
"11010111011100111010010111001110",
"01001110100110111001010000000111",
"11010111011100111010010110000000",
"01001110100110111001010000000111",
"11010111011100111010010111001110",
"11010111011100111010010110000000",
"11101101110001111110101111001110",
"11111011110100000111111001101101",
"11111011110100000111111001101101",
"11111011110100000111111001101101",
"11101101110001111110101111001110",
"11111011110100000111111001101101",
"00001110100001000111101000001011",
"10010100110011110111100110001110",
"10010100110011110111000101000110",
"10010100110011110111100110001110",
"00001110100001000111101000001011",
"10010100110011110111000101000110",
"00000010000001101110000111010100",
"01111100111111111001011110111101",
"01111100111111111001011110111101",
"01111100111111111001011110111101",
"00000010000001101110000111010100",
"01111100111111111001011110111101",
"00110010000100101100110110010101",
"00110100101011111000001001000010",
"00110100101101000001100010101111",
"00110100101011111000001001000010",
"00110010000100101100110110010101",
"00110100101101000001100010101111",
"00100100101011010000001111111001",
"00101110011010111010100010111100",
"00101110011010111010100011010010",
"00101110011010111010100010111100",
"00100100101011010000001111111001",
"00101110011010111010100011010010",
"01000010000001000111100101000101",
"01000000011110100000100000110111",
"01000010000101000001100111001000",
"01000000011110100000100000110111",
"01000010000001000111100101000101",
"01000010000101000001100111001000",
"00101101111101011000010101001100",
"00110010110110100001111111100110",
"00110010110110100101110101000111",
"00110010110110100001111111100110",
"00101101111101011000010101001100",
"00110010110110100101110101000111",
"00101001101010100010111010111110",
"10110100011101000001000100100010",
"10110100011101000001000100011101",
"10110100011101000001000100100010",
"00101001101010100010111010111110",
"10110100011101000001000100011101",
"01011110011101110001010111001011",
"01011100010100000001111101100101",
"01011110100000100000101111100001",
"01011100010100000001111101100101",
"01011110011101110001010111001011",
"01011110100000100000101111100001",
"01110110010001111111111010011011",
"11101010011110000110010011010101",
"01110110010001111111111010011010",
"11101010011110000110010011010101",
"01110110010001111111111010011011",
"01110110010001111111111010011010",
"00110011011010010111001001001101",
"00101110000100111110000110011101",
"00110011011010011001011101000101",
"00101110000100111110000110011101",
"00110011011010010111001001001101",
"00110011011010011001011101000101",
"10110100101000101111001001000111",
"10101110101000010000010110000100",
"10110100101000101111110001010111",
"10101110101000010000010110000100",
"10110100101000101111001001000111",
"10110100101000101111110001010111",
"11110011111110010011101110100101",
"00000001011010101101111101010111",
"11110011111110010011101110100101",
"00000001011010101101111101010111",
"11110011111110010011101110100101",
"11110011111110010011101110100101",
"01100001010110011100101011010001",
"01011011010001111111000101001100",
"01100001010110011101011101010000",
"01011011010001111111000101001100",
"01100001010110011100101011010001",
"01100001010110011101011101010000",
"11010110000101100110111101110000",
"01001011001101100011100000100001",
"11010110000101100110111101101101",
"01001011001101100011100000100001",
"11010110000101100110111101110000",
"11010110000101100110111101101101",
"11001000011100110111110011010000",
"11010111111110111110011101000001",
"11010111111110111110011101000001",
"11010111111110111110011101000001",
"11001000011100110111110011010000",
"11010111111110111110011101000001",
"10000011011000111100001110110110",
"11111001001001011011101011110110",
"11111001001001011011101011110110",
"11111001001001011011101011110110",
"10000011011000111100001110110110",
"11111001001001011011101011110110",
"11100010101111010011110010101100",
"01100111010111100010110100111110",
"01100111010111011100111010100000",
"01100111010111100010110100111110",
"11100010101111010011110010101100",
"01100111010111011100111010100000",
"10010000001001111100000001010001",
"10010100011101001101011010100101",
"10010100011101010111111001100101",
"10010100011101001101011010100101",
"10010000001001111100000001010001",
"10010100011101010111111001100101",
"00011101110001010011111110101010",
"10101010010011100101000100001011",
"10101010010011100101000100001011",
"10101010010011100101000100001011",
"00011101110001010011111110101010",
"10101010010011100101000100001011",
"11110010011110101011001010101000",
"11111001011101101111101100100010",
"11111001011101101111111100001101",
"11111001011101101111101100100010",
"11110010011110101011001010101000",
"11111001011101101111111100001101",
"00011010000111111110111110001001",
"00011011110101111111000110010000",
"00011011111010111110111110000001",
"00011011110101111111000110010000",
"00011010000111111110111110001001",
"00011011111010111110111110000001",
"11000010100100011111000111010000",
"01001010000101110010110110101100",
"01001010000101110010110010001000",
"01001010000101110010110110101100",
"11000010100100011111000111010000",
"01001010000101110010110010001000",
"10100100010100010010001101011111",
"10101110100000110101100101110100",
"10101110100000110101100101111011",
"10101110100000110101100101110100",
"10100100010100010010001101011111",
"10101110100000110101100101111011",
"10100010111000011101010110011101",
"10101110100001110101000101000101",
"10101110100001110101000101000110",
"10101110100001110101000101000101",
"10100010111000011101010110011101",
"10101110100001110101000101000110",
"00110000100010101101111111000001",
"10100001011010111010100101110000",
"00110000100010101101111111000001",
"10100001011010111010100101110000",
"00110000100010101101111111000001",
"00110000100010101101111111000001",
"10110110011110010100111101110010",
"11000101111010111111101010101011",
"11000101111010111111101010101011",
"11000101111010111111101010101011",
"10110110011110010100111101110010",
"11000101111010111111101010101011",
"10100110100110001000100011001001",
"10100111111001100100000110110111",
"10101000000001100011000111110101",
"10100111111001100100000110110111",
"10100110100110001000100011001001",
"10101000000001100011000111110101",
"00010011010101001001100010110110",
"00010110011010001000010011010101",
"00010110011010111101011100111000",
"00010110011010001000010011010101",
"00010011010101001001100010110110",
"00010110011010111101011100111000",
"01110110111001000011110100101111",
"11111100110000101000101001101101",
"11111100110000100111110000101001",
"11111100110000101000101001101101",
"01110110111001000011110100101111",
"11111100110000100111110000101001",
"00110001110100101110100000100101",
"00110111000010001010011001110101",
"00110111000010001100000011010010",
"00110111000010001010011001110101",
"00110001110100101110100000100101",
"00110111000010001100000011010010",
"10001100010011110110001111101110",
"00010111011110100010000110000010",
"00010111011110100010000101111111",
"00010111011110100010000110000010",
"10001100010011110110001111101110",
"00010111011110100010000101111111",
"11011100001100100001010000100000",
"01011001000101010100110001011011",
"11011100001011111011111011101111",
"01011001000101010100110001011011",
"11011100001100100001010000100000",
"11011100001011111011111011101111",
"11001101011010100101101000001110",
"11010100001101011100010010010111",
"11010100001101011100100001000000",
"11010100001101011100010010010111",
"11001101011010100101101000001110",
"11010100001101011100100001000000",
"00010000101111110000010100110010",
"10001101000110101001011100000001",
"00010000101111011101000000000100");

  signal op1,op2,ans1,ans,answ,low,high: std_logic_vector(31 downto 0);
  signal addr: std_logic_vector(9 downto 0) := (others=>'0');
  signal miss: std_logic_vector(31 downto 0) := (others=>'0');
  signal rom_o: std_logic_vector(7 downto 0) := (others=>'1');
  signal uart_go: std_logic;
  signal uart_busy: std_logic := '0';
  signal iter: std_logic_vector(31 downto 0) := (others=>'0');
  signal state: std_logic_vector(4 downto 0) := (others=>'0');
  signal state2: std_logic_vector(4 downto 0) := (others=>'0');

begin

  ib: IBUFG port map (
   i=>MCLK1,
   o=>iclk);
  bg: BUFG port map (
    i=>iclk,
    o=>clk);

  fadder:fadd port map
    (clk, op1, op2, ans);

  rs232c: u232c generic map (wtime=>x"1ADB")
  port map (
    clk=>clk,
    data=>rom_o,
    go=>uart_go,
    busy=>uart_busy,
    tx=>rs_tx);


 cal: process(clk)
 begin
   if rising_edge(clk) then-- hoge clk後に返答
     if state = "00000" then
       state<=state+1;
       addr<=addr+3;
       op1<=rom(conv_integer(addr));
       op2<=rom(conv_integer(addr+1));
       ans1<=rom(conv_integer(addr+2));
     elsif state = "00001" then
       state<=state+1;
     elsif state = "00010" then
       state<=state+1;
       answ<=ans;
       state2<="00000";
     elsif state = "00011" and uart_go = '1'then --op1の出力
       state2<=state2+1;
       if op1(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "00100" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "00101" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "00110" and uart_go = '1'then --op2の出力
       state2<=state2+1;
       if op2(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "00111" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01000" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01001" and uart_go = '1'then --outputの出力
       state2<=state2+1;
       if answ(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01010" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01011" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01100" and uart_go = '1'then --answerの出力
       state2<=state2+1;
       if ans1(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "01101" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "01110" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "01111" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10000" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10001" then --low,highとの比較
       state<=state+1;
       low<=ans1 - 2;
     elsif state = "10010" then
       state<=state+1;
       high<=ans1 + 2;
     elsif state = "10011" then
       iter<=iter+1;
       state<=state+1;
       if high < answ or low > answ then
         miss<=miss+1;
       end if;
     elsif state = "10100" and uart_go = '1'then --iterの出力
       state2<=state2+1;
       if iter(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "10101" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "10110" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "10111" and uart_go = '1'then --missの出力
       state2<=state2+1;
       if miss(31-conv_integer(state2)) = '1' then
         rom_o<=x"31";
       else
         rom_o<=x"30";
       end if;
       if state2 = "11111" then
         state<=state+1;
         state2<="00000";
       end if;
     elsif state = "11000" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11001" and uart_go = '1'then
       state<=state+1;
       rom_o<=x"0a";
     elsif state = "11010" and uart_go = '1'then -- 改行
       state<=state+1;
       rom_o<=x"0d";
     elsif state = "11011" and uart_go = '1'then
       state<="00000";
       rom_o<=x"0a";
     end if;
   end if;
 end process;

    send_msg: process(clk)
  begin
    if rising_edge(clk) then
      if uart_busy='0' and uart_go='0' then
        uart_go<='1';
      else
        uart_go<='0';
      end if;
    end if;
  end process;
  
end VHDL;
