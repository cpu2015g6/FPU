/home/mizuta1018/HW/FPU/VHDL/finv/invromfetch.vhd