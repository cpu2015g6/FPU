library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

entity blockram1 is

  generic (
    dwidth : integer := 23;
    awidth : integer := );

  port (
    clk  : in  std_logic;
    we   : in  std_logic;
    di   : in  std_logic_vector(dwidth - 1 downto 0);
    do   : out std_logic_vector(dwidth - 1 downto 0);
    addr : in  std_logic_vector(awidth - 1 downto 0));

end blockram1;

architecture behavioral of blockram1 is

  type ram_type is
    array(0 to (2 ** awidth) - 1) of std_logic_vector(dwidth - 1 downto 0);

  signal ram : ram_type := (
"01101010000010011110101",
"01101010011001000110000",
"01101010101111101100001",
"01101011000110010000101",
"01101011011100110011111",
"01101011110011010101110",
"01101100001001110110010",
"01101100100000010101010",
"01101100110110110011000",
"01101101001101001111001",
"01101101100011101010001",
"01101101111010000011101",
"01101110010000011011111",
"01101110100110110010100",
"01101110111101001000000",
"01101111010011011100000",
"01101111101001101110110",
"01110000000000000000001",
"01110000010110010000010",
"01110000101100011110111",
"01110001000010101100010",
"01110001011000111000010",
"01110001101111000010111",
"01110010000101001100010",
"01110010011011010100011",
"01110010110001011011001",
"01110011000111100000011",
"01110011011101100100100",
"01110011110011100111001",
"01110100001001101000101",
"01110100011111101000111",
"01110100110101100111110",
"01110101001011100101010",
"01110101100001100001100",
"01110101110111011100100",
"01110110001101010110010",
"01110110100011001110101",
"01110110111001000101101",
"01110111001110111011101",
"01110111100100110000001",
"01110111111010100011100",
"01111000010000010101100",
"01111000100110000110100",
"01111000111011110110001",
"01111001010001100100011",
"01111001100111010001011",
"01111001111100111101001",
"01111010010010100111110",
"01111010101000010001000",
"01111010111101111001001",
"01111011010011011111111",
"01111011101001000101101",
"01111011111110101001111",
"01111100010100001101001",
"01111100101001101111000",
"01111100111111001111111",
"01111101010100101111010",
"01111101101010001101101",
"01111101111111101010101",
"01111110010101000110101",
"01111110101010100001010",
"01111110111111111010110",
"01111111010101010011001",
"01111111101010101010010",
"10000000000000000000010",
"10000000010101010101000",
"10000000101010101000011",
"10000000111111111010110",
"10000001010101001100000",
"10000001101010011100001",
"10000001111111101011000",
"10000010010100111000101",
"10000010101010000101001",
"10000010111111010000101",
"10000011010100011010110",
"10000011101001100011111",
"10000011111110101011110",
"10000100010011110010100",
"10000100101000111000000",
"10000100111101111100100",
"10000101010010111111110",
"10000101101000000010000",
"10000101111101000011001",
"10000110010010000011001",
"10000110100111000001111",
"10000110111011111111100",
"10000111010000111100001",
"10000111100101110111100",
"10000111111010110001110",
"10001000001111101010111",
"10001000100100100011000",
"10001000111001011010000",
"10001001001110001111111",
"10001001100011000100101",
"10001001110111111000010",
"10001010001100101010110",
"10001010100001011100010",
"10001010110110001100110",
"10001011001010111100000",
"10001011011111101010001",
"10001011110100010111010",
"10001100001001000011010",
"10001100011101101110001",
"10001100110010011000001",
"10001101000111000000111",
"10001101011011101000101",
"10001101110000001111010",
"10001110000100110100111",
"10001110011001011001011",
"10001110101101111100111",
"10001111000010011111010",
"10001111010111000000100",
"10001111101011100001000",
"10010000000000000000001",
"10010000010100011110011",
"10010000101000111011100",
"10010000111101010111101",
"10010001010001110010110",
"10010001100110001100110",
"10010001111010100101110",
"10010010001110111101101",
"10010010100011010100110",
"10010010110111101010100",
"10010011001011111111010",
"10010011100000010011001",
"10010011110100100110000",
"10010100001000110111110",
"10010100011101001000101",
"10010100110001011000011",
"10010101000101100111001",
"10010101011001110100111",
"10010101101110000001101",
"10010110000010001101100",
"10010110010110011000001",
"10010110101010100001111",
"10010110111110101010100",
"10010111010010110010011",
"10010111100110111001001",
"10010111111010111110111",
"10011000001111000011101",
"10011000100011000111011",
"10011000110111001010001",
"10011001001011001100000",
"10011001011111001100110",
"10011001110011001100110",
"10011010000111001011110",
"10011010011011001001100",
"10011010101111000110100",
"10011011000011000010100",
"10011011010110111101100",
"10011011101010110111100",
"10011011111110110000101",
"10011100010010101000110",
"10011100100110011111111",
"10011100111010010110001",
"10011101001110001011011",
"10011101100001111111110",
"10011101110101110011000",
"10011110001001100101011",
"10011110011101010110111",
"10011110110001000111100",
"10011111000100110111001",
"10011111011000100101101",
"10011111101100010011011",
"10100000000000000000001",
"10100000010011101100000",
"10100000100111010110111",
"10100000111011000000111",
"10100001001110101010000",
"10100001100010010010000",
"10100001110101111001010",
"10100010001001011111100",
"10100010011101000100111",
"10100010110000101001011",
"10100011000100001100111",
"10100011010111101111100",
"10100011101011010001010",
"10100011111110110010010",
"10100100010010010010001",
"10100100100101110001001",
"10100100111001001111001",
"10100101001100101100011",
"10100101100000001000101",
"10100101110011100100001",
"10100110000110111110101",
"10100110011010011000001",
"10100110101101110000111",
"10100111000001001000110",
"10100111010100011111101",
"10100111100111110101110",
"10100111111011001011000",
"10101000001110011111010",
"10101000100001110010111",
"10101000110101000101010",
"10101001001000010110111",
"10101001011011100111101",
"10101001101110110111110",
"10101010000010000110110",
"10101010010101010101000",
"10101010101000100010010",
"10101010111011101110110",
"10101011001110111010010",
"10101011100010000101001",
"10101011110101001111000",
"10101100001000011000000",
"10101100011011100000001",
"10101100101110100111011",
"10101101000001101101111",
"10101101010100110011100",
"10101101100111111000010",
"10101101111010111100010",
"10101110001101111111010",
"10101110100001000001100",
"10101110110100000010111",
"10101111000111000011101",
"10101111011010000011010",
"10101111101101000010001",
"10110000000000000000001",
"10110000010010111101011",
"10110000100101111001110",
"10110000111000110101010",
"10110001001011110000000",
"10110001011110101010000",
"10110001110001100011000",
"10110010000100011011010",
"10110010010111010010101",
"10110010101010001001010",
"10110010111100111111000",
"10110011001111110100001",
"10110011100010101000010",
"10110011110101011011101",
"10110100001000001110001",
"10110100011010111111111",
"10110100101101110000110",
"10110101000000100001000",
"10110101010011010000010",
"10110101100101111110110",
"10110101111000101100100",
"10110110001011011001011",
"10110110011110000101101",
"10110110110000110000111",
"10110111000011011011011",
"10110111010110000101001",
"10110111101000101110001",
"10110111111011010110001",
"10111000001101111101101",
"10111000100000100100001",
"10111000110011001001111",
"10111001000101101110111",
"10111001011000010011001",
"10111001101010110110101",
"10111001111101011001010",
"10111010001111111011001",
"10111010100010011100010",
"10111010110100111100101",
"10111011000111011100010",
"10111011011001111011001",
"10111011101100011001000",
"10111011111110110110010",
"10111100010001010010111",
"10111100100011101110101",
"10111100110110001001100",
"10111101001000100011110",
"10111101011010111101001",
"10111101101101010101110",
"10111101111111101101110",
"10111110010010000100111",
"10111110100100011011011",
"10111110110110110001000",
"10111111001001000101111",
"10111111011011011010000",
"10111111101101101101100",
"11000000000000000000001",
"11000000010010010010000",
"11000000100100100011001",
"11000000110110110011110",
"11000001001001000011011",
"11000001011011010010011",
"11000001101101100000100",
"11000001111111101101111",
"11000010010001111010101",
"11000010100100000110101",
"11000010110110010001111",
"11000011001000011100100",
"11000011011010100110010",
"11000011101100101111010",
"11000011111110110111101",
"11000100010000111111010",
"11000100100011000110001",
"11000100110101001100010",
"11000101000111010001110",
"11000101011001010110011",
"11000101101011011010011",
"11000101111101011101110",
"11000110001111100000010",
"11000110100001100010001",
"11000110110011100011010",
"11000111000101100011110",
"11000111010111100011011",
"11000111101001100010011",
"11000111111011100000101",
"11001000001101011110010",
"11001000011111011011001",
"11001000110001010111010",
"11001001000011010010110",
"11001001010101001101100",
"11001001100111000111100",
"11001001111001000000111",
"11001010001010111001101",
"11001010011100110001100",
"11001010101110101000110",
"11001011000000011111011",
"11001011010010010101010",
"11001011100100001010011",
"11001011110101111110111",
"11001100000111110010101",
"11001100011001100101110",
"11001100101011011000010",
"11001100111101001010000",
"11001101001110111011000",
"11001101100000101011100",
"11001101110010011011000",
"11001110000100001010001",
"11001110010101111000011",
"11001110100111100110000",
"11001110111001010011000",
"11001111001010111111010",
"11001111011100101010111",
"11001111101110010101111",
"11010000000000000000001",
"11010000010001101001110",
"11010000100011010010101",
"11010000110100111010111",
"11010001000110100010100",
"11010001011000001001011",
"11010001101001101111101",
"11010001111011010101010",
"11010010001100111010001",
"11010010011110011110011",
"11010010110000000010000",
"11010011000001100101000",
"11010011010011000111010",
"11010011100100101001000",
"11010011110110001001111",
"11010100000111101010001",
"11010100011001001001111",
"11010100101010101000111",
"11010100111100000111010",
"11010101001101100100111",
"11010101011111000001111",
"11010101110000011110011",
"11010110000001111010001",
"11010110010011010101010",
"11010110100100101111110",
"11010110110110001001100",
"11010111000111100010110",
"11010111011000111011010",
"11010111101010010011010",
"11010111111011101010011",
"11011000001101000001000",
"11011000011110010111000",
"11011000101111101100011",
"11011001000001000001000",
"11011001010010010101001",
"11011001100011101000101",
"11011001110100111011011",
"11011010000110001101100",
"11011010010111011111001",
"11011010101000110000001",
"11011010111010000000011",
"11011011001011010000001",
"11011011011100011111000",
"11011011101101101101100",
"11011011111110111011010",
"11011100010000001000100",
"11011100100001010101000",
"11011100110010100000111",
"11011101000011101100010",
"11011101010100110110111",
"11011101100110000001000",
"11011101110111001010100",
"11011110001000010011010",
"11011110011001011011100",
"11011110101010100011001",
"11011110111011101010001",
"11011111001100110000100",
"11011111011101110110011",
"11011111101110111011100",
"11100000000000000000001",
"11100000010001000100000",
"11100000100010000111011",
"11100000110011001010001",
"11100001000100001100011",
"11100001010101001110000",
"11100001100110001110110",
"11100001110111001111000",
"11100010001000001111000",
"11100010011001001110000",
"11100010101010001100101",
"11100010111011001010101",
"11100011001100001000000",
"11100011011101000100101",
"11100011101110000000111",
"11100011111110111100011",
"11100100001111110111011",
"11100100100000110001110",
"11100100110001101011100",
"11100101000010100100110",
"11100101010011011101011",
"11100101100100010101011",
"11100101110101001100111",
"11100110000110000011110",
"11100110010110111010000",
"11100110100111101111110",
"11100110111000100100111",
"11100111001001011001011",
"11100111011010001101011",
"11100111101011000000110",
"11100111111011110011100",
"11101000001100100101110",
"11101000011101010111011",
"11101000101110001000011",
"11101000111110111000110",
"11101001001111101000111",
"11101001100000011000010",
"11101001110001000111000",
"11101010000001110101001",
"11101010010010100010110",
"11101010100011001111110",
"11101010110011111100010",
"11101011000100101000010",
"11101011010101010011101",
"11101011100101111110011",
"11101011110110101000101",
"11101100000111010010010",
"11101100010111111011011",
"11101100101000100011111",
"11101100111001001011111",
"11101101001001110011010",
"11101101011010011010001",
"11101101101011000000011",
"11101101111011100110001",
"11101110001100001011011",
"11101110011100110000000",
"11101110101101010100000",
"11101110111101110111100",
"11101111001110011010100",
"11101111011110111100111",
"11101111101111011110110",
"11110000000000000000001",
"11110000010000100000111",
"11110000100001000001001",
"11110000110001100000110",
"11110001000001111111111",
"11110001010010011110100",
"11110001100010111100100",
"11110001110011011001111",
"11110010000011110110111",
"11110010010100010011010",
"11110010100100101111000",
"11110010110101001010011",
"11110011000101100101001",
"11110011010101111111011",
"11110011100110011001000",
"11110011110110110010001",
"11110100000111001010110",
"11110100010111100010111",
"11110100100111111010011",
"11110100111000010001011",
"11110101001000100111111",
"11110101011000111101110",
"11110101101001010011010",
"11110101111001101000001",
"11110110001001111100011",
"11110110011010010000010",
"11110110101010100011100",
"11110110111010110110010",
"11110111001011001000101",
"11110111011011011010010",
"11110111101011101011011",
"11110111111011111100000",
"11111000001100001100001",
"11111000011100011011110",
"11111000101100101010111",
"11111000111100111001011",
"11111001001101000111011",
"11111001011101010100111",
"11111001101101100001111",
"11111001111101101110011",
"11111010001101111010011",
"11111010011110000101110",
"11111010101110010000110",
"11111010111110011011001",
"11111011001110100101000",
"11111011011110101110011",
"11111011101110110111010",
"11111011111110111111101",
"11111100001111000111011",
"11111100011111001110110",
"11111100101111010101101",
"11111100111111011011111",
"11111101001111100001101",
"11111101011111100111000",
"11111101101111101011110",
"11111101111111110000000",
"11111110001111110011110",
"11111110011111110111001",
"11111110101111111001111",
"11111110111111111100001",
"11111111001111111101111",
"11111111011111111111001",
"11111111101111111111111",
"00000000000000000000000",
"00000000001111111111101",
"00000000011111111110001",
"00000000101111111011101",
"00000000111111111000001",
"00000001001111110011101",
"00000001011111101110010",
"00000001101111100111110",
"00000001111111100000011",
"00000010001111011000000",
"00000010011111001110101",
"00000010101111000100010",
"00000010111110111001000",
"00000011001110101100101",
"00000011011110011111011",
"00000011101110010001010",
"00000011111110000010000",
"00000100001101110010000",
"00000100011101100000111",
"00000100101101001110111",
"00000100111100111011111",
"00000101001100101000000",
"00000101011100010011001",
"00000101101011111101011",
"00000101111011100110101",
"00000110001011001110111",
"00000110011010110110100",
"00000110101010011101000",
"00000110111010000010100",
"00000111001001100111001",
"00000111011001001010111",
"00000111101000101101101",
"00000111111000001111100",
"00001000000111110000100",
"00001000010111010000101",
"00001000100110101111101",
"00001000110110001101111",
"00001001000101101011010",
"00001001010101000111110",
"00001001100100100011010",
"00001001110011111101111",
"00001010000011010111101",
"00001010010010110000100",
"00001010100010001000101",
"00001010110001011111101",
"00001011000000110101111",
"00001011010000001011001",
"00001011011111011111101",
"00001011101110110011001",
"00001011111110000101111",
"00001100001101010111101",
"00001100011100101000101",
"00001100101011111000110",
"00001100111011000111111",
"00001101001010010110010",
"00001101011001100011110",
"00001101101000110000011",
"00001101110111111100001",
"00001110000111000111001",
"00001110010110010001010",
"00001110100101011010011",
"00001110110100100010110",
"00001111000011101010011",
"00001111010010110001000",
"00001111100001110110111",
"00001111110000111100000",
"00010000000000000000001",
"00010000001111000011100",
"00010000011110000110000",
"00010000101101000111101",
"00010000111100001000100",
"00010001001011001000100",
"00010001011010000111110",
"00010001101001000110010",
"00010001111000000011110",
"00010010000111000000100",
"00010010010101111100011",
"00010010100100110111100",
"00010010110011110001111",
"00010011000010101011011",
"00010011010001100100001",
"00010011100000011100000",
"00010011101111010011001",
"00010011111110001001011",
"00010100001100111110111",
"00010100011011110011100",
"00010100101010100111100",
"00010100111001011010101",
"00010101001000001100111",
"00010101010110111110100",
"00010101100101101111010",
"00010101110100011111010",
"00010110000011001110011",
"00010110010001111100110",
"00010110100000101010011",
"00010110101111010111010",
"00010110111110000011011",
"00010111001100101110101",
"00010111011011011001001",
"00010111101010000010111",
"00010111111000101011111",
"00011000000111010100001",
"00011000010101111011101",
"00011000100100100010010",
"00011000110011001000010",
"00011001000001101101011",
"00011001010000010001111",
"00011001011110110101100",
"00011001101101011000100",
"00011001111011111010101",
"00011010001010011100000",
"00011010011000111100110",
"00011010100111011100110",
"00011010110101111011111",
"00011011000100011010010",
"00011011010010111000000",
"00011011100001010101000",
"00011011101111110001010",
"00011011111110001100110",
"00011100001100100111100",
"00011100011011000001100",
"00011100101001011010110",
"00011100110111110011011",
"00011101000110001011010",
"00011101010100100010011",
"00011101100010111000110",
"00011101110001001110100",
"00011101111111100011011",
"00011110001101110111110",
"00011110011100001011010",
"00011110101010011110000",
"00011110111000110000001",
"00011111000111000001101",
"00011111010101010010010",
"00011111100011100010010",
"00011111110001110001100",
"00100000000000000000001",
"00100000001110001110000",
"00100000011100011011001",
"00100000101010100111101",
"00100000111000110011011",
"00100001000110111110100",
"00100001010101001000111",
"00100001100011010010100",
"00100001110001011011100",
"00100001111111100011111",
"00100010001101101011100",
"00100010011011110010011",
"00100010101001111000101",
"00100010110111111110010",
"00100011000110000011001",
"00100011010100000111010",
"00100011100010001010111",
"00100011110000001101110",
"00100011111110001111111",
"00100100001100010001011",
"00100100011010010010010",
"00100100101000010010011",
"00100100110110010001111",
"00100101000100010000101",
"00100101010010001110111",
"00100101100000001100010",
"00100101101110001001001",
"00100101111100000101010",
"00100110001010000000110",
"00100110010111111011101",
"00100110100101110101111",
"00100110110011101111011",
"00100111000001101000010",
"00100111001111100000100",
"00100111011101011000000",
"00100111101011001110111",
"00100111111001000101010",
"00101000000110111010111",
"00101000010100101111110",
"00101000100010100100001",
"00101000110000010111111",
"00101000111110001010111",
"00101001001011111101010",
"00101001011001101111000",
"00101001100111100000001",
"00101001110101010000101",
"00101010000011000000100",
"00101010010000101111110",
"00101010011110011110011",
"00101010101100001100010",
"00101010111001111001101",
"00101011000111100110010",
"00101011010101010010011",
"00101011100010111101111",
"00101011110000101000101",
"00101011111110010010111",
"00101100001011111100011",
"00101100011001100101011",
"00101100100111001101110",
"00101100110100110101100",
"00101101000010011100101",
"00101101010000000011001",
"00101101011101101001000",
"00101101101011001110010",
"00101101111000110010111",
"00101110000110010110111",
"00101110010011111010011",
"00101110100001011101001",
"00101110101110111111011",
"00101110111100100001000",
"00101111001010000010000",
"00101111010111100010100",
"00101111100101000010010",
"00101111110010100001100",
"00110000000000000000001",
"00110000001101011110001",
"00110000011010111011100",
"00110000101000011000011",
"00110000110101110100101",
"00110001000011010000010",
"00110001010000101011010",
"00110001011110000101110",
"00110001101011011111101",
"00110001111000111000111",
"00110010000110010001101",
"00110010010011101001110",
"00110010100001000001010",
"00110010101110011000001",
"00110010111011101110100",
"00110011001001000100011",
"00110011010110011001100",
"00110011100011101110001",
"00110011110001000010010",
"00110011111110010101110",
"00110100001011101000101",
"00110100011000111010111",
"00110100100110001100101",
"00110100110011011101111",
"00110101000000101110100",
"00110101001101111110100",
"00110101011011001110000",
"00110101101000011100111",
"00110101110101101011010",
"00110110000010111001000",
"00110110010000000110010",
"00110110011101010010111",
"00110110101010011111000",
"00110110110111101010101",
"00110111000100110101100",
"00110111010010000000000",
"00110111011111001001111",
"00110111101100010011001",
"00110111111001011011111",
"00111000000110100100001",
"00111000010011101011110",
"00111000100000110010111",
"00111000101101111001011",
"00111000111010111111011",
"00111001001000000100111",
"00111001010101001001110",
"00111001100010001110001",
"00111001101111010010000",
"00111001111100010101010",
"00111010001001011000000",
"00111010010110011010010",
"00111010100011011011111",
"00111010110000011101000",
"00111010111101011101100",
"00111011001010011101101",
"00111011010111011101001",
"00111011100100011100000",
"00111011110001011010100",
"00111011111110011000011",
"00111100001011010101110",
"00111100011000010010101",
"00111100100101001110111",
"00111100110010001010110",
"00111100111111000110000",
"00111101001100000000101",
"00111101011000111010111",
"00111101100101110100100",
"00111101110010101101110",
"00111101111111100110011",
"00111110001100011110011",
"00111110011001010110000",
"00111110100110001101001",
"00111110110011000011101",
"00111110111111111001101",
"00111111001100101111001",
"00111111011001100100001",
"00111111100110011000101",
"00111111110011001100101",
"01000000000000000000001",
"01000000001100110011000",
"01000000011001100101100",
"01000000100110010111011",
"01000000110011001000110",
"01000000111111111001110",
"01000001001100101010001",
"01000001011001011010000",
"01000001100110001001011",
"01000001110010111000001",
"01000001111111100110101",
"01000010001100010100100",
"01000010011001000001111",
"01000010100101101110110",
"01000010110010011011001",
"01000010111111000111000",
"01000011001011110010011",
"01000011011000011101010",
"01000011100101000111101",
"01000011110001110001100",
"01000011111110011011000",
"01000100001011000011111",
"01000100010111101100010",
"01000100100100010100001",
"01000100110000111011101",
"01000100111101100010100",
"01000101001010001001000",
"01000101010110101111000",
"01000101100011010100011",
"01000101101111111001011",
"01000101111100011101111",
"01000110001001000001111",
"01000110010101100101100",
"01000110100010001000100",
"01000110101110101011001",
"01000110111011001101001",
"01000111000111101110110",
"01000111010100001111111",
"01000111100000110000100",
"01000111101101010000110",
"01000111111001110000011",
"01001000000110001111101",
"01001000010010101110011",
"01001000011111001100101",
"01001000101011101010100",
"01001000111000000111110",
"01001001000100100100101",
"01001001010001000001000",
"01001001011101011100111",
"01001001101001111000011",
"01001001110110010011011",
"01001010000010101101111",
"01001010001111000111111",
"01001010011011100001100",
"01001010100111111010101",
"01001010110100010011010",
"01001011000000101011011",
"01001011001101000011001",
"01001011011001011010011",
"01001011100101110001001",
"01001011110010000111100",
"01001011111110011101011",
"01001100001010110010110",
"01001100010111000111110",
"01001100100011011100010",
"01001100101111110000011",
"01001100111100000011111",
"01001101001000010111000",
"01001101010100101001110",
"01001101100000111100000",
"01001101101101001101110",
"01001101111001011111001",
"01001110000101110000000",
"01001110010010000000011",
"01001110011110010000011",
"01001110101010011111111",
"01001110110110101111000",
"01001111000010111101101",
"01001111001111001011110",
"01001111011011011001100",
"01001111100111100110110",
"01001111110011110011101",
"01010000000000000000001",
"01010000001100001100000",
"01010000011000010111101",
"01010000100100100010101",
"01010000110000101101011",
"01010000111100110111100",
"01010001001001000001010",
"01010001010101001010101",
"01010001100001010011100",
"01010001101101011100000",
"01010001111001100100000",
"01010010000101101011101",
"01010010010001110010110",
"01010010011101111001100",
"01010010101001111111110",
"01010010110110000101101",
"01010011000010001011000",
"01010011001110010000000",
"01010011011010010100101",
"01010011100110011000110",
"01010011110010011100011",
"01010011111110011111110",
"01010100001010100010100",
"01010100010110100101000",
"01010100100010100111000",
"01010100101110101000100",
"01010100111010101001110",
"01010101000110101010011",
"01010101010010101010110",
"01010101011110101010101",
"01010101101010101010001",
"01010101110110101001001",
"01010110000010100111110",
"01010110001110100110000",
"01010110011010100011110",
"01010110100110100001001",
"01010110110010011110000",
"01010110111110011010101",
"01010111001010010110110",
"01010111010110010010011",
"01010111100010001101101",
"01010111101110001000100",
"01010111111010000011000",
"01011000000101111101000",
"01011000010001110110110",
"01011000011101101111111",
"01011000101001101000110",
"01011000110101100001001",
"01011001000001011001001",
"01011001001101010000110",
"01011001011001000111111",
"01011001100100111110101",
"01011001110000110101000",
"01011001111100101011000",
"01011010001000100000100",
"01011010010100010101101",
"01011010100000001010011",
"01011010101011111110110",
"01011010110111110010110",
"01011011000011100110010",
"01011011001111011001011",
"01011011011011001100001",
"01011011100110111110100",
"01011011110010110000011",
"01011011111110100001111",
"01011100001010010011000",
"01011100010110000011110",
"01011100100001110100001",
"01011100101101100100001",
"01011100111001010011101",
"01011101000101000010110",
"01011101010000110001100",
"01011101011100011111111",
"01011101101000001101111",
"01011101110011111011100",
"01011101111111101000101",
"01011110001011010101100",
"01011110010111000001111",
"01011110100010101101111",
"01011110101110011001100",
"01011110111010000100110",
"01011111000101101111100",
"01011111010001011010001",
"01011111011101000100001",
"01011111101000101101111",
"01011111110100010111001",
"01100000000000000000000",
"01100000001011101000101",
"01100000010111010000110",
"01100000100010111000100",
"01100000101110011111111",
"01100000111010000110111",
"01100001000101101101100",
"01100001010001010011110",
"01100001011100111001101",
"01100001101000011111001",
"01100001110100000100010",
"01100001111111101001000",
"01100010001011001101010",
"01100010010110110001010",
"01100010100010010100111",
"01100010101101111000000",
"01100010111001011010111",
"01100011000100111101011",
"01100011010000011111011",
"01100011011100000001001",
"01100011100111100010100",
"01100011110011000011100",
"01100011111110100100000",
"01100100001010000100010",
"01100100010101100100001",
"01100100100001000011101",
"01100100101100100010110",
"01100100111000000001011",
"01100101000011011111110",
"01100101001110111101110",
"01100101011010011011011",
"01100101100101111000110",
"01100101110001010101101",
"01100101111100110010001",
"01100110001000001110010",
"01100110010011101010001",
"01100110011111000101100",
"01100110101010100000101",
"01100110110101111011010",
"01100111000001010101101",
"01100111001100101111101",
"01100111011000001001010",
"01100111100011100010100",
"01100111101110111011011",
"01100111111010010100000",
"01101000000101101100001",
"01101000010001000100000",
"01101000011100011011011",
"01101000100111110010100",
"01101000110011001001010",
"01101000111110011111101",
"01101001001001110101101",
"01101001010101001011011",
"01101001100000100000101",
"01101001101011110101101",
"01101001110111001010010");

  signal reg_addr : std_logic_vector(awidth - 1 downto 0);

begin

  process(clk)
  begin
    if rising_edge(clk) then
      if we = '1' then
        ram(conv_integer(addr)) <= di;
      end if;
      reg_addr <= addr;
    end if;
  end process;

  do <= ram(conv_integer(reg_addr));

end behavioral;
